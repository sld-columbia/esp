../../cores/ariane/ariane/src/common_cells/src/sram.sv