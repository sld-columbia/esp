fasdf
