-- AMBA Wrapper for Xilinx System Monitor
  constant CFG_GRSYSMON : integer := CONFIG_GRSYSMON;

