-- Xilinx MIG
  constant CFG_MIG_DDR2    : integer := CONFIG_MIG_DDR2;
  constant CFG_MIG_RANKS   : integer := CONFIG_MIG_RANKS;
  constant CFG_MIG_COLBITS : integer := CONFIG_MIG_COLBITS;
  constant CFG_MIG_ROWBITS : integer := CONFIG_MIG_ROWBITS;
  constant CFG_MIG_BANKBITS: integer := CONFIG_MIG_BANKBITS;
  constant CFG_MIG_HMASK   : integer := 16#CONFIG_MIG_HMASK#;


