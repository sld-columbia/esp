#include "grlib_config.h"
#include "tkconfig.h"

  -----------------------------------------------------------------------------
  --  LEON3 Demonstration design test bench configuration
  --  Copyright (C) 2009 Aeroflex Gaisler
  ------------------------------------------------------------------------------
  use work.gencomp.all;

package grlib_config is

#include "grlib_config.vhd.h"

end package grlib_config;
