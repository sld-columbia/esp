../ariane/ariane/src/register_interface/src/reg_intf_pkg.sv