`ifndef VX_FPU_DEFINE
`define VX_FPU_DEFINE

`include "VX_define.vh"

`IGNORE_WARNINGS_BEGIN
import fpu_types::*;
`IGNORE_WARNINGS_END

`endif
