../vortex/hw/rtl/cache/VX_cache_define.vh