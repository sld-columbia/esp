../vortex/hw/rtl/VX_define.vh