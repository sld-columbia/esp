
library ieee;
use ieee.std_logic_1164.all;
library unisim;
use unisim.vcomponents.all;

entity virtex4_mul_61x61 is
port(
  A : in std_logic_vector(60 downto 0);
  B : in std_logic_vector(60 downto 0);
  EN :  in std_logic;
  CLK :  in std_logic;
  PRODUCT : out std_logic_vector(121 downto 0));
end virtex4_mul_61x61;

architecture beh of virtex4_mul_61x61 is
  signal R1IN_3_2_1 : std_logic_vector(33 downto 17);
  signal R1IN_3_2 : std_logic_vector(16 downto 0);
  signal R1IN_2_2_1 : std_logic_vector(33 downto 17);
  signal R1IN_2_2 : std_logic_vector(16 downto 0);
  signal R1IN_4_4_2 : std_logic_vector(26 downto 0);
  signal R1IN_ADD_1 : std_logic_vector(31 downto 0);
  signal R1IN_4 : std_logic_vector(52 downto 17);
  signal R1IN_4_3_1 : std_logic_vector(33 downto 17);
  signal R1IN_4_3 : std_logic_vector(16 downto 0);
  signal R1IN_4_2 : std_logic_vector(16 downto 0);
  signal R1IN_4_2_1 : std_logic_vector(33 downto 17);
  signal R1IN_4_2F : std_logic_vector(43 downto 1);
  signal R1IN_4_3F : std_logic_vector(43 downto 0);
  signal R1IN_1FF : std_logic_vector(33 downto 18);
  signal R1IN_4FF : std_logic_vector(16 downto 0);
  signal R1IN_2_2F : std_logic_vector(43 downto 1);
  signal R1IN_4_4_ADD_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_4_4_ADD_1_PCOUT : std_logic_vector(47 downto 0);
  signal R1IN_2_2_ADD_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_2_2_ADD_1_PCOUT : std_logic_vector(47 downto 0);
  signal R1IN_3_2_ADD_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_3_2_ADD_1_PCOUT : std_logic_vector(47 downto 0);
  signal R1IN_4_2_ADD_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_4_2_ADD_1_PCOUT : std_logic_vector(47 downto 0);
  signal R1IN_4_3_ADD_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_4_3_ADD_1_PCOUT : std_logic_vector(47 downto 0);
  signal R1IN_4_4_2_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_2_2_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_3_2_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_4_2_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_4_3_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_1_PCOUT : std_logic_vector(47 downto 0);
  signal R1IN_2_1_PCOUT : std_logic_vector(47 downto 0);
  signal R1IN_3_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_3_1_PCOUT : std_logic_vector(47 downto 0);
  signal R1IN_4_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_4_1_PCOUT : std_logic_vector(47 downto 0);
  signal R1IN_4_4_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_4_4_1_PCOUT : std_logic_vector(47 downto 0);
  signal R1IN_4_4_4_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_4_4_4_PCOUT : std_logic_vector(47 downto 0);
  signal R1IN_4_4_2_0 : std_logic_vector(26 downto 0);
  signal R1IN_2_2_0 : std_logic_vector(16 downto 0);
  signal R1IN_2_2_1_0 : std_logic_vector(33 downto 17);
  signal R1IN_3_2_0 : std_logic_vector(16 downto 0);
  signal R1IN_3_2_1_0 : std_logic_vector(33 downto 17);
  signal R1IN_4_2_0 : std_logic_vector(16 downto 0);
  signal R1IN_4_2_1_0 : std_logic_vector(33 downto 17);
  signal R1IN_4_3_0 : std_logic_vector(16 downto 0);
  signal R1IN_4_3_1_0 : std_logic_vector(33 downto 17);
  signal B_0 : std_logic_vector(16 downto 0);
  signal R1IN_4_4 : std_logic_vector(53 downto 17);
  signal R1IN_2F_RETO : std_logic_vector(16 downto 0);
  signal R1IN_3F : std_logic_vector(16 downto 0);
  signal R1IN_3F_RETO : std_logic_vector(16 downto 0);
  signal R1IN_2_RETO : std_logic_vector(60 downto 17);
  signal R1IN_3_1F_RETO : std_logic_vector(33 downto 17);
  signal R1IN_3 : std_logic_vector(60 downto 17);
  signal R1IN_4_1F_RETO : std_logic_vector(33 downto 17);
  signal R1IN_4_ADD_1_RETO : std_logic_vector(44 downto 1);
  signal R1IN_4_4F : std_logic_vector(16 downto 0);
  signal R1IN_4_4F_RETO : std_logic_vector(16 downto 0);
  signal R1IN_4_4_ADD_1F_RETO : std_logic_vector(27 downto 0);
  signal R1IN_3_1F : std_logic_vector(33 downto 17);
  signal R1IN_3_1F_RETO_0 : std_logic_vector(17 to 17);
  signal R1IN_3_2F : std_logic_vector(43 downto 1);
  signal R1IN_3_2F_RETO : std_logic_vector(43 downto 1);
  signal R1IN_4_4_ADD_1F : std_logic_vector(27 downto 0);
  signal R1IN_4_4_ADD_1F_RETO_0 : std_logic_vector(0 to 0);
  signal R1IN_4_4_1F : std_logic_vector(33 downto 18);
  signal R1IN_4_4_1F_RETO : std_logic_vector(33 downto 18);
  signal R1IN_4_4_4F_RETO : std_logic_vector(19 downto 0);
  signal R1IN_4_4_4_P : std_logic_vector(47 downto 20);
  signal R1IN_4_1_P : std_logic_vector(47 downto 34);
  signal R1IN_2_1F_RETO : std_logic_vector(33 downto 17);
  signal R1IN_2_2F_RETO : std_logic_vector(43 downto 1);
  signal R1IN_4_3F_RETO : std_logic_vector(43 downto 0);
  signal R1IN_4_2F_RETO : std_logic_vector(43 downto 1);
  signal R1IN_2_1_P : std_logic_vector(47 downto 34);
  signal NN_1 : std_logic ;
  signal NN_2 : std_logic ;
  signal R1IN_4_ADD_1 : std_logic ;
  signal R1IN_ADD_2 : std_logic ;
  signal R1IN_2_ADD_1 : std_logic ;
  signal UC : std_logic ;
  signal UC_0 : std_logic ;
  signal UC_1 : std_logic ;
  signal UC_2 : std_logic ;
  signal UC_3 : std_logic ;
  signal UC_4 : std_logic ;
  signal UC_5 : std_logic ;
  signal UC_6 : std_logic ;
  signal UC_7 : std_logic ;
  signal UC_8 : std_logic ;
  signal UC_9 : std_logic ;
  signal UC_10 : std_logic ;
  signal UC_11 : std_logic ;
  signal UC_12 : std_logic ;
  signal UC_13 : std_logic ;
  signal UC_14 : std_logic ;
  signal UC_15 : std_logic ;
  signal UC_16 : std_logic ;
  signal UC_17 : std_logic ;
  signal UC_18 : std_logic ;
  signal UC_19 : std_logic ;
  signal UC_20 : std_logic ;
  signal UC_21 : std_logic ;
  signal UC_22 : std_logic ;
  signal UC_23 : std_logic ;
  signal UC_24 : std_logic ;
  signal UC_25 : std_logic ;
  signal UC_26 : std_logic ;
  signal UC_27 : std_logic ;
  signal UC_28 : std_logic ;
  signal UC_29 : std_logic ;
  signal UC_30 : std_logic ;
  signal UC_31 : std_logic ;
  signal UC_32 : std_logic ;
  signal UC_33 : std_logic ;
  signal UC_34 : std_logic ;
  signal UC_35 : std_logic ;
  signal UC_36 : std_logic ;
  signal UC_37 : std_logic ;
  signal UC_38 : std_logic ;
  signal UC_39 : std_logic ;
  signal UC_40 : std_logic ;
  signal UC_41 : std_logic ;
  signal UC_42 : std_logic ;
  signal UC_43 : std_logic ;
  signal UC_44 : std_logic ;
  signal UC_45 : std_logic ;
  signal UC_46 : std_logic ;
  signal UC_47 : std_logic ;
  signal UC_48 : std_logic ;
  signal UC_49 : std_logic ;
  signal UC_50 : std_logic ;
  signal UC_51 : std_logic ;
  signal UC_52 : std_logic ;
  signal UC_53 : std_logic ;
  signal UC_54 : std_logic ;
  signal UC_55 : std_logic ;
  signal UC_56 : std_logic ;
  signal UC_57 : std_logic ;
  signal UC_58 : std_logic ;
  signal UC_59 : std_logic ;
  signal UC_60 : std_logic ;
  signal UC_61 : std_logic ;
  signal UC_62 : std_logic ;
  signal UC_63 : std_logic ;
  signal UC_64 : std_logic ;
  signal UC_65 : std_logic ;
  signal UC_66 : std_logic ;
  signal UC_67 : std_logic ;
  signal UC_68 : std_logic ;
  signal UC_69 : std_logic ;
  signal UC_70 : std_logic ;
  signal UC_71 : std_logic ;
  signal UC_72 : std_logic ;
  signal UC_73 : std_logic ;
  signal UC_74 : std_logic ;
  signal UC_75 : std_logic ;
  signal UC_76 : std_logic ;
  signal UC_77 : std_logic ;
  signal UC_78 : std_logic ;
  signal UC_79 : std_logic ;
  signal UC_80 : std_logic ;
  signal UC_81 : std_logic ;
  signal UC_82 : std_logic ;
  signal UC_83 : std_logic ;
  signal UC_84 : std_logic ;
  signal UC_85 : std_logic ;
  signal UC_86 : std_logic ;
  signal UC_87 : std_logic ;
  signal UC_88 : std_logic ;
  signal UC_89 : std_logic ;
  signal UC_90 : std_logic ;
  signal UC_91 : std_logic ;
  signal UC_92 : std_logic ;
  signal UC_93 : std_logic ;
  signal UC_94 : std_logic ;
  signal UC_95 : std_logic ;
  signal UC_96 : std_logic ;
  signal UC_97 : std_logic ;
  signal UC_98 : std_logic ;
  signal UC_99 : std_logic ;
  signal UC_100 : std_logic ;
  signal UC_101 : std_logic ;
  signal UC_102 : std_logic ;
  signal UC_103 : std_logic ;
  signal UC_104 : std_logic ;
  signal UC_105 : std_logic ;
  signal UC_106 : std_logic ;
  signal UC_107 : std_logic ;
  signal UC_108 : std_logic ;
  signal UC_109 : std_logic ;
  signal UC_110 : std_logic ;
  signal UC_111 : std_logic ;
  signal UC_112 : std_logic ;
  signal UC_113 : std_logic ;
  signal UC_114 : std_logic ;
  signal UC_115 : std_logic ;
  signal UC_116 : std_logic ;
  signal UC_117 : std_logic ;
  signal UC_118 : std_logic ;
  signal UC_119 : std_logic ;
  signal UC_120 : std_logic ;
  signal UC_121 : std_logic ;
  signal UC_122 : std_logic ;
  signal UC_123 : std_logic ;
  signal UC_124 : std_logic ;
  signal UC_125 : std_logic ;
  signal UC_126 : std_logic ;
  signal UC_127 : std_logic ;
  signal UC_128 : std_logic ;
  signal UC_129 : std_logic ;
  signal UC_130 : std_logic ;
  signal UC_131 : std_logic ;
  signal UC_132 : std_logic ;
  signal UC_133 : std_logic ;
  signal UC_134 : std_logic ;
  signal UC_135 : std_logic ;
  signal UC_136 : std_logic ;
  signal UC_137 : std_logic ;
  signal UC_138 : std_logic ;
  signal UC_139 : std_logic ;
  signal UC_140 : std_logic ;
  signal UC_141 : std_logic ;
  signal UC_142 : std_logic ;
  signal UC_143 : std_logic ;
  signal UC_144 : std_logic ;
  signal UC_145 : std_logic ;
  signal UC_146 : std_logic ;
  signal UC_147 : std_logic ;
  signal UC_148 : std_logic ;
  signal UC_149 : std_logic ;
  signal UC_150 : std_logic ;
  signal UC_151 : std_logic ;
  signal UC_152 : std_logic ;
  signal UC_153 : std_logic ;
  signal UC_154 : std_logic ;
  signal UC_155 : std_logic ;
  signal UC_156 : std_logic ;
  signal UC_157 : std_logic ;
  signal UC_158 : std_logic ;
  signal UC_159 : std_logic ;
  signal UC_160 : std_logic ;
  signal UC_161 : std_logic ;
  signal UC_162 : std_logic ;
  signal UC_163 : std_logic ;
  signal UC_164 : std_logic ;
  signal UC_165 : std_logic ;
  signal UC_166 : std_logic ;
  signal UC_167 : std_logic ;
  signal UC_168 : std_logic ;
  signal UC_169 : std_logic ;
  signal UC_170 : std_logic ;
  signal UC_171 : std_logic ;
  signal UC_172 : std_logic ;
  signal UC_173 : std_logic ;
  signal UC_174 : std_logic ;
  signal UC_175 : std_logic ;
  signal UC_176 : std_logic ;
  signal UC_177 : std_logic ;
  signal UC_178 : std_logic ;
  signal UC_179 : std_logic ;
  signal UC_180 : std_logic ;
  signal UC_181 : std_logic ;
  signal UC_182 : std_logic ;
  signal UC_183 : std_logic ;
  signal UC_184 : std_logic ;
  signal UC_185 : std_logic ;
  signal UC_186 : std_logic ;
  signal UC_187 : std_logic ;
  signal UC_188 : std_logic ;
  signal UC_189 : std_logic ;
  signal UC_190 : std_logic ;
  signal UC_191 : std_logic ;
  signal UC_192 : std_logic ;
  signal UC_193 : std_logic ;
  signal UC_208 : std_logic ;
  signal UC_209 : std_logic ;
  signal UC_210 : std_logic ;
  signal UC_211 : std_logic ;
  signal UC_212 : std_logic ;
  signal UC_213 : std_logic ;
  signal UC_214 : std_logic ;
  signal UC_215 : std_logic ;
  signal UC_216 : std_logic ;
  signal UC_217 : std_logic ;
  signal UC_218 : std_logic ;
  signal UC_219 : std_logic ;
  signal UC_220 : std_logic ;
  signal UC_221 : std_logic ;
  signal UC_236 : std_logic ;
  signal UC_237 : std_logic ;
  signal UC_238 : std_logic ;
  signal UC_239 : std_logic ;
  signal UC_240 : std_logic ;
  signal UC_241 : std_logic ;
  signal UC_242 : std_logic ;
  signal UC_243 : std_logic ;
  signal UC_244 : std_logic ;
  signal UC_245 : std_logic ;
  signal UC_246 : std_logic ;
  signal UC_247 : std_logic ;
  signal UC_248 : std_logic ;
  signal UC_249 : std_logic ;
  signal UC_103_0 : std_logic ;
  signal UC_104_0 : std_logic ;
  signal UC_105_0 : std_logic ;
  signal UC_106_0 : std_logic ;
  signal UC_107_0 : std_logic ;
  signal UC_108_0 : std_logic ;
  signal UC_109_0 : std_logic ;
  signal UC_110_0 : std_logic ;
  signal UC_111_0 : std_logic ;
  signal UC_112_0 : std_logic ;
  signal UC_113_0 : std_logic ;
  signal UC_114_0 : std_logic ;
  signal UC_115_0 : std_logic ;
  signal UC_116_0 : std_logic ;
  signal UC_117_0 : std_logic ;
  signal UC_118_0 : std_logic ;
  signal UC_119_0 : std_logic ;
  signal UC_120_0 : std_logic ;
  signal UC_121_0 : std_logic ;
  signal UC_122_0 : std_logic ;
  signal UC_123_0 : std_logic ;
  signal UC_124_0 : std_logic ;
  signal UC_125_0 : std_logic ;
  signal UC_126_0 : std_logic ;
  signal UC_127_0 : std_logic ;
  signal UC_128_0 : std_logic ;
  signal UC_129_0 : std_logic ;
  signal UC_130_0 : std_logic ;
  signal UC_131_0 : std_logic ;
  signal UC_132_0 : std_logic ;
  signal UC_133_0 : std_logic ;
  signal UC_134_0 : std_logic ;
  signal UC_135_0 : std_logic ;
  signal UC_136_0 : std_logic ;
  signal UC_137_0 : std_logic ;
  signal UC_138_0 : std_logic ;
  signal UC_139_0 : std_logic ;
  signal UC_140_0 : std_logic ;
  signal UC_141_0 : std_logic ;
  signal UC_142_0 : std_logic ;
  signal UC_143_0 : std_logic ;
  signal UC_144_0 : std_logic ;
  signal UC_145_0 : std_logic ;
  signal UC_146_0 : std_logic ;
  signal UC_147_0 : std_logic ;
  signal UC_148_0 : std_logic ;
  signal UC_149_0 : std_logic ;
  signal UC_150_0 : std_logic ;
  signal UC_151_0 : std_logic ;
  signal UC_152_0 : std_logic ;
  signal UC_153_0 : std_logic ;
  signal UC_154_0 : std_logic ;
  signal UC_155_0 : std_logic ;
  signal UC_156_0 : std_logic ;
  signal UC_157_0 : std_logic ;
  signal UC_158_0 : std_logic ;
  signal UC_159_0 : std_logic ;
  signal UC_160_0 : std_logic ;
  signal UC_161_0 : std_logic ;
  signal UC_162_0 : std_logic ;
  signal UC_163_0 : std_logic ;
  signal UC_164_0 : std_logic ;
  signal UC_165_0 : std_logic ;
  signal UC_166_0 : std_logic ;
  signal UC_167_0 : std_logic ;
  signal UC_168_0 : std_logic ;
  signal UC_169_0 : std_logic ;
  signal UC_170_0 : std_logic ;
  signal UC_171_0 : std_logic ;
  signal UC_172_0 : std_logic ;
  signal UC_173_0 : std_logic ;
  signal UC_174_0 : std_logic ;
  signal UC_175_0 : std_logic ;
  signal UC_176_0 : std_logic ;
  signal UC_177_0 : std_logic ;
  signal UC_178_0 : std_logic ;
  signal UC_179_0 : std_logic ;
  signal GND_0 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_0 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_1 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_1 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_2 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_2 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_3 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_3 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_4 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_4 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_5 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_5 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_6 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_6 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_7 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_7 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_8 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_8 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_9 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_9 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_10 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_10 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_11 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_11 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_12 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_12 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_13 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_13 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_14 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_14 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_15 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_15 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_16 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_16 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_17 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_17 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_18 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_18 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_19 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_19 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_20 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_20 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_21 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_21 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_22 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_22 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_23 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_23 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_24 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_24 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_25 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_25 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_26 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_26 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_27 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_27 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_28 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_28 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_29 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_29 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_30 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_30 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_31 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_31 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_32 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_32 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_33 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_33 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_34 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_34 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_35 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_0 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_1 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_1 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_2 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_2 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_3 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_3 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_4 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_4 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_5 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_5 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_6 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_6 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_7 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_7 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_8 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_8 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_9 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_9 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_10 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_10 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_11 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_11 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_12 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_12 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_13 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_13 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_14 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_14 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_15 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_15 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_16 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_16 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_17 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_17 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_18 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_18 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_19 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_19 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_20 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_20 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_21 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_21 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_22 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_22 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_23 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_23 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_24 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_24 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_25 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_25 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_26 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_26 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_27 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_27 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_28 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_28 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_29 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_29 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_30 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_30 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_31 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_31 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_32 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_32 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_33 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_33 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_34 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_0 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_1 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_1 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_2 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_2 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_3 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_3 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_4 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_4 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_5 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_5 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_6 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_6 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_7 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_7 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_8 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_8 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_9 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_9 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_10 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_10 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_11 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_11 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_12 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_12 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_13 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_13 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_14 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_14 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_15 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_15 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_16 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_16 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_17 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_17 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_18 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_18 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_19 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_19 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_20 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_20 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_21 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_21 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_22 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_22 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_23 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_23 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_24 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_24 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_25 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_25 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_26 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_26 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_27 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_27 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_28 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_28 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_29 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_29 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_30 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_30 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_31 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_31 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_32 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_32 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_33 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_33 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_34 : std_logic ;
  signal R1IN_ADD_1_0_CRY_0 : std_logic ;
  signal R1IN_ADD_1_0_AXB_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_1 : std_logic ;
  signal R1IN_ADD_1_0_AXB_2 : std_logic ;
  signal R1IN_ADD_1_0_CRY_2 : std_logic ;
  signal R1IN_ADD_1_0_AXB_3 : std_logic ;
  signal R1IN_ADD_1_0_CRY_3 : std_logic ;
  signal R1IN_ADD_1_0_AXB_4 : std_logic ;
  signal R1IN_ADD_1_0_CRY_4 : std_logic ;
  signal R1IN_ADD_1_0_AXB_5 : std_logic ;
  signal R1IN_ADD_1_0_CRY_5 : std_logic ;
  signal R1IN_ADD_1_0_AXB_6 : std_logic ;
  signal R1IN_ADD_1_0_CRY_6 : std_logic ;
  signal R1IN_ADD_1_0_AXB_7 : std_logic ;
  signal R1IN_ADD_1_0_CRY_7 : std_logic ;
  signal R1IN_ADD_1_0_AXB_8 : std_logic ;
  signal R1IN_ADD_1_0_CRY_8 : std_logic ;
  signal R1IN_ADD_1_0_AXB_9 : std_logic ;
  signal R1IN_ADD_1_0_CRY_9 : std_logic ;
  signal R1IN_ADD_1_0_AXB_10 : std_logic ;
  signal R1IN_ADD_1_0_CRY_10 : std_logic ;
  signal R1IN_ADD_1_0_AXB_11 : std_logic ;
  signal R1IN_ADD_1_0_CRY_11 : std_logic ;
  signal R1IN_ADD_1_0_AXB_12 : std_logic ;
  signal R1IN_ADD_1_0_CRY_12 : std_logic ;
  signal R1IN_ADD_1_0_AXB_13 : std_logic ;
  signal R1IN_ADD_1_0_CRY_13 : std_logic ;
  signal R1IN_ADD_1_0_AXB_14 : std_logic ;
  signal R1IN_ADD_1_0_CRY_14 : std_logic ;
  signal R1IN_ADD_1_0_AXB_15 : std_logic ;
  signal R1IN_ADD_1_0_CRY_15 : std_logic ;
  signal R1IN_ADD_1_0_AXB_16 : std_logic ;
  signal R1IN_ADD_1_0_CRY_16 : std_logic ;
  signal R1IN_ADD_1_0_AXB_17 : std_logic ;
  signal R1IN_ADD_1_0_CRY_17 : std_logic ;
  signal R1IN_ADD_1_0_AXB_18 : std_logic ;
  signal R1IN_ADD_1_0_CRY_18 : std_logic ;
  signal R1IN_ADD_1_0_AXB_19 : std_logic ;
  signal R1IN_ADD_1_0_CRY_19 : std_logic ;
  signal R1IN_ADD_1_0_AXB_20 : std_logic ;
  signal R1IN_ADD_1_0_CRY_20 : std_logic ;
  signal R1IN_ADD_1_0_AXB_21 : std_logic ;
  signal R1IN_ADD_1_0_CRY_21 : std_logic ;
  signal R1IN_ADD_1_0_AXB_22 : std_logic ;
  signal R1IN_ADD_1_0_CRY_22 : std_logic ;
  signal R1IN_ADD_1_0_AXB_23 : std_logic ;
  signal R1IN_ADD_1_0_CRY_23 : std_logic ;
  signal R1IN_ADD_1_0_AXB_24 : std_logic ;
  signal R1IN_ADD_1_0_CRY_24 : std_logic ;
  signal R1IN_ADD_1_0_AXB_25 : std_logic ;
  signal R1IN_ADD_1_0_CRY_25 : std_logic ;
  signal R1IN_ADD_1_0_AXB_26 : std_logic ;
  signal R1IN_ADD_1_0_CRY_26 : std_logic ;
  signal R1IN_ADD_1_0_AXB_27 : std_logic ;
  signal R1IN_ADD_1_0_CRY_27 : std_logic ;
  signal R1IN_ADD_1_0_AXB_28 : std_logic ;
  signal R1IN_ADD_1_0_CRY_28 : std_logic ;
  signal R1IN_ADD_1_0_AXB_29 : std_logic ;
  signal R1IN_ADD_1_0_CRY_29 : std_logic ;
  signal R1IN_ADD_1_0_AXB_30 : std_logic ;
  signal R1IN_ADD_1_0_CRY_30 : std_logic ;
  signal R1IN_ADD_1_0_AXB_31 : std_logic ;
  signal R1IN_ADD_1_1_CRY_0 : std_logic ;
  signal R1IN_ADD_1_1_AXB_1 : std_logic ;
  signal R1IN_ADD_1_1_CRY_1 : std_logic ;
  signal R1IN_ADD_1_1_AXB_2 : std_logic ;
  signal R1IN_ADD_1_1_CRY_2 : std_logic ;
  signal R1IN_ADD_1_1_AXB_3 : std_logic ;
  signal R1IN_ADD_1_1_CRY_3 : std_logic ;
  signal R1IN_ADD_1_1_AXB_4 : std_logic ;
  signal R1IN_ADD_1_1_CRY_4 : std_logic ;
  signal R1IN_ADD_1_1_AXB_5 : std_logic ;
  signal R1IN_ADD_1_1_CRY_5 : std_logic ;
  signal R1IN_ADD_1_1_AXB_6 : std_logic ;
  signal R1IN_ADD_1_1_CRY_6 : std_logic ;
  signal R1IN_ADD_1_1_AXB_7 : std_logic ;
  signal R1IN_ADD_1_1_CRY_7 : std_logic ;
  signal R1IN_ADD_1_1_AXB_8 : std_logic ;
  signal R1IN_ADD_1_1_CRY_8 : std_logic ;
  signal R1IN_ADD_1_1_AXB_9 : std_logic ;
  signal R1IN_ADD_1_1_CRY_9 : std_logic ;
  signal R1IN_ADD_1_1_AXB_10 : std_logic ;
  signal R1IN_ADD_1_1_CRY_10 : std_logic ;
  signal R1IN_ADD_1_1_AXB_11 : std_logic ;
  signal R1IN_ADD_1_1_CRY_11 : std_logic ;
  signal R1IN_ADD_1_1_AXB_12 : std_logic ;
  signal R1IN_ADD_1_1_CRY_12 : std_logic ;
  signal R1IN_ADD_1_1_AXB_13 : std_logic ;
  signal R1IN_ADD_1_1_CRY_13 : std_logic ;
  signal R1IN_ADD_1_1_AXB_14 : std_logic ;
  signal R1IN_ADD_1_1_CRY_14 : std_logic ;
  signal R1IN_ADD_1_1_AXB_15 : std_logic ;
  signal R1IN_ADD_1_1_CRY_15 : std_logic ;
  signal R1IN_ADD_1_1_AXB_16 : std_logic ;
  signal R1IN_ADD_1_1_CRY_16 : std_logic ;
  signal R1IN_ADD_1_1_AXB_17 : std_logic ;
  signal R1IN_ADD_1_1_CRY_17 : std_logic ;
  signal R1IN_ADD_1_1_AXB_18 : std_logic ;
  signal R1IN_ADD_1_1_CRY_18 : std_logic ;
  signal R1IN_ADD_1_1_AXB_19 : std_logic ;
  signal R1IN_ADD_1_1_CRY_19 : std_logic ;
  signal R1IN_ADD_1_1_AXB_20 : std_logic ;
  signal R1IN_ADD_1_1_CRY_20 : std_logic ;
  signal R1IN_ADD_1_1_AXB_21 : std_logic ;
  signal R1IN_ADD_1_1_CRY_21 : std_logic ;
  signal R1IN_ADD_1_1_AXB_22 : std_logic ;
  signal R1IN_ADD_1_1_CRY_22 : std_logic ;
  signal R1IN_ADD_1_1_AXB_23 : std_logic ;
  signal R1IN_ADD_1_1_CRY_23 : std_logic ;
  signal R1IN_ADD_1_1_AXB_24 : std_logic ;
  signal R1IN_ADD_1_1_CRY_24 : std_logic ;
  signal R1IN_ADD_1_1_AXB_25 : std_logic ;
  signal R1IN_ADD_1_1_CRY_25 : std_logic ;
  signal R1IN_ADD_1_1_AXB_26 : std_logic ;
  signal R1IN_ADD_1_1_CRY_26 : std_logic ;
  signal R1IN_ADD_1_1_AXB_27 : std_logic ;
  signal R1IN_ADD_1_1_CRY_27 : std_logic ;
  signal R1IN_ADD_1_1_AXB_28 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_0 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_1 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_1 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_2 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_2 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_3 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_3 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_4 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_4 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_5 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_5 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_6 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_6 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_7 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_7 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_8 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_8 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_9 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_9 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_10 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_10 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_11 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_11 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_12 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_12 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_13 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_13 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_14 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_14 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_15 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_15 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_16 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_16 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_17 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_17 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_18 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_18 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_19 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_19 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_20 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_20 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_21 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_21 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_22 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_22 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_23 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_23 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_24 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_24 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_25 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_25 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_26 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_26 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_27 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_27 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_28 : std_logic ;
  signal R1IN_3_ADD_1_CRY_0 : std_logic ;
  signal R1IN_3_ADD_1_AXB_1 : std_logic ;
  signal R1IN_3_ADD_1_CRY_1 : std_logic ;
  signal R1IN_3_ADD_1_AXB_2 : std_logic ;
  signal R1IN_3_ADD_1_CRY_2 : std_logic ;
  signal R1IN_3_ADD_1_AXB_3 : std_logic ;
  signal R1IN_3_ADD_1_CRY_3 : std_logic ;
  signal R1IN_3_ADD_1_AXB_4 : std_logic ;
  signal R1IN_3_ADD_1_CRY_4 : std_logic ;
  signal R1IN_3_ADD_1_AXB_5 : std_logic ;
  signal R1IN_3_ADD_1_CRY_5 : std_logic ;
  signal R1IN_3_ADD_1_AXB_6 : std_logic ;
  signal R1IN_3_ADD_1_CRY_6 : std_logic ;
  signal R1IN_3_ADD_1_AXB_7 : std_logic ;
  signal R1IN_3_ADD_1_CRY_7 : std_logic ;
  signal R1IN_3_ADD_1_AXB_8 : std_logic ;
  signal R1IN_3_ADD_1_CRY_8 : std_logic ;
  signal R1IN_3_ADD_1_AXB_9 : std_logic ;
  signal R1IN_3_ADD_1_CRY_9 : std_logic ;
  signal R1IN_3_ADD_1_AXB_10 : std_logic ;
  signal R1IN_3_ADD_1_CRY_10 : std_logic ;
  signal R1IN_3_ADD_1_AXB_11 : std_logic ;
  signal R1IN_3_ADD_1_CRY_11 : std_logic ;
  signal R1IN_3_ADD_1_AXB_12 : std_logic ;
  signal R1IN_3_ADD_1_CRY_12 : std_logic ;
  signal R1IN_3_ADD_1_AXB_13 : std_logic ;
  signal R1IN_3_ADD_1_CRY_13 : std_logic ;
  signal R1IN_3_ADD_1_AXB_14 : std_logic ;
  signal R1IN_3_ADD_1_CRY_14 : std_logic ;
  signal R1IN_3_ADD_1_AXB_15 : std_logic ;
  signal R1IN_3_ADD_1_CRY_15 : std_logic ;
  signal R1IN_3_ADD_1_AXB_16 : std_logic ;
  signal R1IN_3_ADD_1_CRY_16 : std_logic ;
  signal R1IN_3_ADD_1_AXB_17 : std_logic ;
  signal R1IN_3_ADD_1_CRY_17 : std_logic ;
  signal R1IN_3_ADD_1_AXB_18 : std_logic ;
  signal R1IN_3_ADD_1_CRY_18 : std_logic ;
  signal R1IN_3_ADD_1_AXB_19 : std_logic ;
  signal R1IN_3_ADD_1_CRY_19 : std_logic ;
  signal R1IN_3_ADD_1_AXB_20 : std_logic ;
  signal R1IN_3_ADD_1_CRY_20 : std_logic ;
  signal R1IN_3_ADD_1_AXB_21 : std_logic ;
  signal R1IN_3_ADD_1_CRY_21 : std_logic ;
  signal R1IN_3_ADD_1_AXB_22 : std_logic ;
  signal R1IN_3_ADD_1_CRY_22 : std_logic ;
  signal R1IN_3_ADD_1_AXB_23 : std_logic ;
  signal R1IN_3_ADD_1_CRY_23 : std_logic ;
  signal R1IN_3_ADD_1_AXB_24 : std_logic ;
  signal R1IN_3_ADD_1_CRY_24 : std_logic ;
  signal R1IN_3_ADD_1_AXB_25 : std_logic ;
  signal R1IN_3_ADD_1_CRY_25 : std_logic ;
  signal R1IN_3_ADD_1_AXB_26 : std_logic ;
  signal R1IN_3_ADD_1_CRY_26 : std_logic ;
  signal R1IN_3_ADD_1_AXB_27 : std_logic ;
  signal R1IN_3_ADD_1_CRY_27 : std_logic ;
  signal R1IN_3_ADD_1_AXB_28 : std_logic ;
  signal R1IN_3_ADD_1_CRY_28 : std_logic ;
  signal R1IN_3_ADD_1_AXB_29 : std_logic ;
  signal R1IN_3_ADD_1_CRY_29 : std_logic ;
  signal R1IN_3_ADD_1_AXB_30 : std_logic ;
  signal R1IN_3_ADD_1_CRY_30 : std_logic ;
  signal R1IN_3_ADD_1_AXB_31 : std_logic ;
  signal R1IN_3_ADD_1_CRY_31 : std_logic ;
  signal R1IN_3_ADD_1_AXB_32 : std_logic ;
  signal R1IN_3_ADD_1_CRY_32 : std_logic ;
  signal R1IN_3_ADD_1_AXB_33 : std_logic ;
  signal R1IN_3_ADD_1_CRY_33 : std_logic ;
  signal R1IN_3_ADD_1_AXB_34 : std_logic ;
  signal R1IN_3_ADD_1_CRY_34 : std_logic ;
  signal R1IN_3_ADD_1_AXB_35 : std_logic ;
  signal R1IN_3_ADD_1_CRY_35 : std_logic ;
  signal R1IN_3_ADD_1_AXB_36 : std_logic ;
  signal R1IN_3_ADD_1_CRY_36 : std_logic ;
  signal R1IN_3_ADD_1_AXB_37 : std_logic ;
  signal R1IN_3_ADD_1_CRY_37 : std_logic ;
  signal R1IN_3_ADD_1_AXB_38 : std_logic ;
  signal R1IN_3_ADD_1_CRY_38 : std_logic ;
  signal R1IN_3_ADD_1_AXB_39 : std_logic ;
  signal R1IN_3_ADD_1_CRY_39 : std_logic ;
  signal R1IN_3_ADD_1_AXB_40 : std_logic ;
  signal R1IN_3_ADD_1_CRY_40 : std_logic ;
  signal R1IN_3_ADD_1_AXB_41 : std_logic ;
  signal R1IN_3_ADD_1_CRY_41 : std_logic ;
  signal R1IN_3_ADD_1_AXB_42 : std_logic ;
  signal R1IN_3_ADD_1_CRY_42 : std_logic ;
  signal R1IN_3_ADD_1_AXB_43 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_0 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_1 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_1 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_2 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_2 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_3 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_3 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_4 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_4 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_5 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_5 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_6 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_6 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_7 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_7 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_8 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_8 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_9 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_9 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_10 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_10 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_11 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_11 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_12 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_12 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_13 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_13 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_14 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_14 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_15 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_15 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_16 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_16 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_17 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_17 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_18 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_18 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_19 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_19 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_20 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_20 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_21 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_21 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_22 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_22 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_23 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_23 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_24 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_24 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_25 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_25 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_26 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_26 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_27 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_27 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_28 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_28 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_29 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_29 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_30 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_30 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_31 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_31 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_32 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_32 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_33 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_33 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_34 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_34 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_35 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_35 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_36 : std_logic ;
  signal NN_3 : std_logic ;
  signal R1IN_ADD_2_CRY_0 : std_logic ;
  signal R1IN_ADD_2_AXB_1 : std_logic ;
  signal R1IN_ADD_2_CRY_1 : std_logic ;
  signal R1IN_ADD_2_AXB_2 : std_logic ;
  signal R1IN_ADD_2_CRY_2 : std_logic ;
  signal R1IN_ADD_2_AXB_3 : std_logic ;
  signal R1IN_ADD_2_CRY_3 : std_logic ;
  signal R1IN_ADD_2_AXB_4 : std_logic ;
  signal R1IN_ADD_2_CRY_4 : std_logic ;
  signal R1IN_ADD_2_AXB_5 : std_logic ;
  signal R1IN_ADD_2_CRY_5 : std_logic ;
  signal R1IN_ADD_2_AXB_6 : std_logic ;
  signal R1IN_ADD_2_CRY_6 : std_logic ;
  signal R1IN_ADD_2_AXB_7 : std_logic ;
  signal R1IN_ADD_2_CRY_7 : std_logic ;
  signal R1IN_ADD_2_AXB_8 : std_logic ;
  signal R1IN_ADD_2_CRY_8 : std_logic ;
  signal R1IN_ADD_2_AXB_9 : std_logic ;
  signal R1IN_ADD_2_CRY_9 : std_logic ;
  signal R1IN_ADD_2_AXB_10 : std_logic ;
  signal R1IN_ADD_2_CRY_10 : std_logic ;
  signal R1IN_ADD_2_AXB_11 : std_logic ;
  signal R1IN_ADD_2_CRY_11 : std_logic ;
  signal R1IN_ADD_2_AXB_12 : std_logic ;
  signal R1IN_ADD_2_CRY_12 : std_logic ;
  signal R1IN_ADD_2_AXB_13 : std_logic ;
  signal R1IN_ADD_2_CRY_13 : std_logic ;
  signal R1IN_ADD_2_AXB_14 : std_logic ;
  signal R1IN_ADD_2_CRY_14 : std_logic ;
  signal R1IN_ADD_2_AXB_15 : std_logic ;
  signal R1IN_ADD_2_CRY_15 : std_logic ;
  signal R1IN_ADD_2_AXB_16 : std_logic ;
  signal R1IN_ADD_2_CRY_16 : std_logic ;
  signal R1IN_ADD_2_AXB_17 : std_logic ;
  signal R1IN_ADD_2_CRY_17 : std_logic ;
  signal R1IN_ADD_2_AXB_18 : std_logic ;
  signal R1IN_ADD_2_CRY_18 : std_logic ;
  signal R1IN_ADD_2_AXB_19 : std_logic ;
  signal R1IN_ADD_2_CRY_19 : std_logic ;
  signal R1IN_ADD_2_AXB_20 : std_logic ;
  signal R1IN_ADD_2_CRY_20 : std_logic ;
  signal R1IN_ADD_2_AXB_21 : std_logic ;
  signal R1IN_ADD_2_CRY_21 : std_logic ;
  signal R1IN_ADD_2_AXB_22 : std_logic ;
  signal R1IN_ADD_2_CRY_22 : std_logic ;
  signal R1IN_ADD_2_AXB_23 : std_logic ;
  signal R1IN_ADD_2_CRY_23 : std_logic ;
  signal R1IN_ADD_2_AXB_24 : std_logic ;
  signal R1IN_ADD_2_CRY_24 : std_logic ;
  signal R1IN_ADD_2_AXB_25 : std_logic ;
  signal R1IN_ADD_2_CRY_25 : std_logic ;
  signal R1IN_ADD_2_AXB_26 : std_logic ;
  signal R1IN_ADD_2_CRY_26 : std_logic ;
  signal R1IN_ADD_2_AXB_27 : std_logic ;
  signal R1IN_ADD_2_CRY_27 : std_logic ;
  signal R1IN_ADD_2_AXB_28 : std_logic ;
  signal R1IN_ADD_2_CRY_28 : std_logic ;
  signal R1IN_ADD_2_AXB_29 : std_logic ;
  signal R1IN_ADD_2_CRY_29 : std_logic ;
  signal R1IN_ADD_2_AXB_30 : std_logic ;
  signal R1IN_ADD_2_CRY_30 : std_logic ;
  signal R1IN_ADD_2_AXB_31 : std_logic ;
  signal R1IN_ADD_2_CRY_31 : std_logic ;
  signal R1IN_ADD_2_AXB_32 : std_logic ;
  signal R1IN_ADD_2_CRY_32 : std_logic ;
  signal R1IN_ADD_2_AXB_33 : std_logic ;
  signal R1IN_ADD_2_CRY_33 : std_logic ;
  signal R1IN_ADD_2_AXB_34 : std_logic ;
  signal R1IN_ADD_2_CRY_34 : std_logic ;
  signal R1IN_ADD_2_AXB_35 : std_logic ;
  signal R1IN_ADD_2_CRY_35 : std_logic ;
  signal R1IN_ADD_2_AXB_36 : std_logic ;
  signal R1IN_ADD_2_CRY_36 : std_logic ;
  signal R1IN_ADD_2_AXB_37 : std_logic ;
  signal R1IN_ADD_2_CRY_37 : std_logic ;
  signal R1IN_ADD_2_AXB_38 : std_logic ;
  signal R1IN_ADD_2_CRY_38 : std_logic ;
  signal R1IN_ADD_2_AXB_39 : std_logic ;
  signal R1IN_ADD_2_CRY_39 : std_logic ;
  signal R1IN_ADD_2_AXB_40 : std_logic ;
  signal R1IN_ADD_2_CRY_40 : std_logic ;
  signal R1IN_ADD_2_AXB_41 : std_logic ;
  signal R1IN_ADD_2_CRY_41 : std_logic ;
  signal R1IN_ADD_2_AXB_42 : std_logic ;
  signal R1IN_ADD_2_CRY_42 : std_logic ;
  signal R1IN_ADD_2_AXB_43 : std_logic ;
  signal R1IN_ADD_2_CRY_43 : std_logic ;
  signal R1IN_ADD_2_AXB_44 : std_logic ;
  signal R1IN_ADD_2_CRY_44 : std_logic ;
  signal R1IN_ADD_2_AXB_45 : std_logic ;
  signal R1IN_ADD_2_CRY_45 : std_logic ;
  signal R1IN_ADD_2_AXB_46 : std_logic ;
  signal R1IN_ADD_2_CRY_46 : std_logic ;
  signal R1IN_ADD_2_AXB_47 : std_logic ;
  signal R1IN_ADD_2_CRY_47 : std_logic ;
  signal R1IN_ADD_2_AXB_48 : std_logic ;
  signal R1IN_ADD_2_CRY_48 : std_logic ;
  signal R1IN_ADD_2_AXB_49 : std_logic ;
  signal R1IN_ADD_2_CRY_49 : std_logic ;
  signal R1IN_ADD_2_AXB_50 : std_logic ;
  signal R1IN_ADD_2_CRY_50 : std_logic ;
  signal R1IN_ADD_2_AXB_51 : std_logic ;
  signal R1IN_ADD_2_CRY_51 : std_logic ;
  signal R1IN_ADD_2_AXB_52 : std_logic ;
  signal R1IN_ADD_2_CRY_52 : std_logic ;
  signal R1IN_ADD_2_AXB_53 : std_logic ;
  signal R1IN_ADD_2_CRY_53 : std_logic ;
  signal R1IN_ADD_2_AXB_54 : std_logic ;
  signal R1IN_ADD_2_CRY_54 : std_logic ;
  signal R1IN_ADD_2_AXB_55 : std_logic ;
  signal R1IN_ADD_2_CRY_55 : std_logic ;
  signal R1IN_ADD_2_AXB_56 : std_logic ;
  signal R1IN_ADD_2_CRY_56 : std_logic ;
  signal R1IN_ADD_2_AXB_57 : std_logic ;
  signal R1IN_ADD_2_CRY_57 : std_logic ;
  signal R1IN_ADD_2_AXB_58 : std_logic ;
  signal R1IN_ADD_2_CRY_58 : std_logic ;
  signal R1IN_ADD_2_AXB_59 : std_logic ;
  signal R1IN_ADD_2_CRY_59 : std_logic ;
  signal R1IN_ADD_2_AXB_60 : std_logic ;
  signal R1IN_ADD_2_CRY_60 : std_logic ;
  signal R1IN_ADD_2_AXB_61 : std_logic ;
  signal R1IN_ADD_2_CRY_61 : std_logic ;
  signal R1IN_ADD_2_AXB_62 : std_logic ;
  signal R1IN_ADD_2_CRY_62 : std_logic ;
  signal R1IN_ADD_2_AXB_63 : std_logic ;
  signal R1IN_ADD_2_CRY_63 : std_logic ;
  signal R1IN_ADD_2_AXB_64 : std_logic ;
  signal R1IN_ADD_2_CRY_64 : std_logic ;
  signal R1IN_ADD_2_AXB_65 : std_logic ;
  signal R1IN_ADD_2_CRY_65 : std_logic ;
  signal R1IN_ADD_2_AXB_66 : std_logic ;
  signal R1IN_ADD_2_CRY_66 : std_logic ;
  signal R1IN_ADD_2_AXB_67 : std_logic ;
  signal R1IN_ADD_2_CRY_67 : std_logic ;
  signal R1IN_ADD_2_AXB_68 : std_logic ;
  signal R1IN_ADD_2_CRY_68 : std_logic ;
  signal R1IN_ADD_2_AXB_69 : std_logic ;
  signal R1IN_ADD_2_CRY_69 : std_logic ;
  signal R1IN_ADD_2_AXB_70 : std_logic ;
  signal R1IN_ADD_2_CRY_70 : std_logic ;
  signal R1IN_ADD_2_AXB_71 : std_logic ;
  signal R1IN_ADD_2_CRY_71 : std_logic ;
  signal R1IN_ADD_2_AXB_72 : std_logic ;
  signal R1IN_ADD_2_CRY_72 : std_logic ;
  signal R1IN_ADD_2_AXB_73 : std_logic ;
  signal R1IN_ADD_2_CRY_73 : std_logic ;
  signal R1IN_ADD_2_AXB_74 : std_logic ;
  signal R1IN_ADD_2_CRY_74 : std_logic ;
  signal R1IN_ADD_2_AXB_75 : std_logic ;
  signal R1IN_ADD_2_CRY_75 : std_logic ;
  signal R1IN_ADD_2_AXB_76 : std_logic ;
  signal R1IN_ADD_2_CRY_76 : std_logic ;
  signal R1IN_ADD_2_AXB_77 : std_logic ;
  signal R1IN_ADD_2_CRY_77 : std_logic ;
  signal R1IN_ADD_2_AXB_78 : std_logic ;
  signal R1IN_ADD_2_CRY_78 : std_logic ;
  signal R1IN_ADD_2_AXB_79 : std_logic ;
  signal R1IN_ADD_2_CRY_79 : std_logic ;
  signal R1IN_ADD_2_AXB_80 : std_logic ;
  signal R1IN_ADD_2_CRY_80 : std_logic ;
  signal R1IN_ADD_2_AXB_81 : std_logic ;
  signal R1IN_ADD_2_CRY_81 : std_logic ;
  signal R1IN_ADD_2_AXB_82 : std_logic ;
  signal R1IN_ADD_2_CRY_82 : std_logic ;
  signal R1IN_ADD_2_AXB_83 : std_logic ;
  signal R1IN_ADD_2_CRY_83 : std_logic ;
  signal R1IN_ADD_2_AXB_84 : std_logic ;
  signal R1IN_ADD_2_CRY_84 : std_logic ;
  signal R1IN_ADD_2_AXB_85 : std_logic ;
  signal R1IN_ADD_2_CRY_85 : std_logic ;
  signal R1IN_ADD_2_AXB_86 : std_logic ;
  signal R1IN_ADD_2_CRY_86 : std_logic ;
  signal R1IN_ADD_2_AXB_87 : std_logic ;
  signal R1IN_ADD_2_CRY_87 : std_logic ;
  signal R1IN_ADD_2_AXB_88 : std_logic ;
  signal R1IN_ADD_2_CRY_88 : std_logic ;
  signal R1IN_ADD_2_AXB_89 : std_logic ;
  signal R1IN_ADD_2_CRY_89 : std_logic ;
  signal R1IN_ADD_2_AXB_90 : std_logic ;
  signal R1IN_ADD_2_CRY_90 : std_logic ;
  signal R1IN_ADD_2_AXB_91 : std_logic ;
  signal R1IN_ADD_2_CRY_91 : std_logic ;
  signal R1IN_ADD_2_AXB_92 : std_logic ;
  signal R1IN_ADD_2_CRY_92 : std_logic ;
  signal R1IN_ADD_2_AXB_93 : std_logic ;
  signal R1IN_ADD_2_CRY_93 : std_logic ;
  signal R1IN_ADD_2_AXB_94 : std_logic ;
  signal R1IN_ADD_2_CRY_94 : std_logic ;
  signal R1IN_ADD_2_AXB_95 : std_logic ;
  signal R1IN_ADD_2_CRY_95 : std_logic ;
  signal R1IN_ADD_2_AXB_96 : std_logic ;
  signal R1IN_ADD_2_CRY_96 : std_logic ;
  signal R1IN_ADD_2_AXB_97 : std_logic ;
  signal R1IN_ADD_2_CRY_97 : std_logic ;
  signal R1IN_ADD_2_AXB_98 : std_logic ;
  signal R1IN_ADD_2_CRY_98 : std_logic ;
  signal R1IN_ADD_2_AXB_99 : std_logic ;
  signal R1IN_ADD_2_CRY_99 : std_logic ;
  signal R1IN_ADD_2_AXB_100 : std_logic ;
  signal R1IN_ADD_2_CRY_100 : std_logic ;
  signal R1IN_ADD_2_AXB_101 : std_logic ;
  signal R1IN_ADD_2_CRY_101 : std_logic ;
  signal R1IN_ADD_2_AXB_102 : std_logic ;
  signal R1IN_ADD_2_CRY_102 : std_logic ;
  signal R1IN_ADD_2_AXB_103 : std_logic ;
  signal R1IN_ADD_2_CRY_103 : std_logic ;
  signal R1IN_ADD_2_AXB_104 : std_logic ;
  signal N_1433 : std_logic ;
  signal N_1592 : std_logic ;
  signal N_4634 : std_logic ;
  signal N_1431 : std_logic ;
  signal N_1591 : std_logic ;
  signal N_4635 : std_logic ;
  signal N_1429 : std_logic ;
  signal N_1590 : std_logic ;
  signal N_4636 : std_logic ;
  signal N_1427 : std_logic ;
  signal N_1589 : std_logic ;
  signal N_4637 : std_logic ;
  signal N_1425 : std_logic ;
  signal N_1588 : std_logic ;
  signal N_4638 : std_logic ;
  signal N_1423 : std_logic ;
  signal N_1587 : std_logic ;
  signal N_4639 : std_logic ;
  signal N_1421 : std_logic ;
  signal N_1586 : std_logic ;
  signal N_4640 : std_logic ;
  signal N_1419 : std_logic ;
  signal N_1585 : std_logic ;
  signal N_4641 : std_logic ;
  signal N_1511 : std_logic ;
  signal N_1556 : std_logic ;
  signal N_4642 : std_logic ;
  signal N_1417 : std_logic ;
  signal N_1584 : std_logic ;
  signal N_4643 : std_logic ;
  signal N_1509 : std_logic ;
  signal N_1555 : std_logic ;
  signal N_4644 : std_logic ;
  signal N_1415 : std_logic ;
  signal N_1583 : std_logic ;
  signal N_4645 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_28 : std_logic ;
  signal R1IN_ADD_1_1_CRY_28 : std_logic ;
  signal N_4646 : std_logic ;
  signal N_1507 : std_logic ;
  signal N_1554 : std_logic ;
  signal N_4647 : std_logic ;
  signal N_1413 : std_logic ;
  signal N_1582 : std_logic ;
  signal N_4648 : std_logic ;
  signal N_1505 : std_logic ;
  signal N_1553 : std_logic ;
  signal N_4649 : std_logic ;
  signal N_1411 : std_logic ;
  signal N_1581 : std_logic ;
  signal N_4650 : std_logic ;
  signal N_1503 : std_logic ;
  signal N_1552 : std_logic ;
  signal N_4651 : std_logic ;
  signal N_1409 : std_logic ;
  signal N_1580 : std_logic ;
  signal N_4652 : std_logic ;
  signal N_1501 : std_logic ;
  signal N_1551 : std_logic ;
  signal N_4653 : std_logic ;
  signal N_1407 : std_logic ;
  signal N_1579 : std_logic ;
  signal N_4654 : std_logic ;
  signal N_1499 : std_logic ;
  signal N_1550 : std_logic ;
  signal N_4655 : std_logic ;
  signal N_1405 : std_logic ;
  signal N_1578 : std_logic ;
  signal N_4656 : std_logic ;
  signal N_1497 : std_logic ;
  signal N_1549 : std_logic ;
  signal N_4657 : std_logic ;
  signal N_1403 : std_logic ;
  signal N_1577 : std_logic ;
  signal N_4658 : std_logic ;
  signal N_1495 : std_logic ;
  signal N_1548 : std_logic ;
  signal N_4659 : std_logic ;
  signal N_1401 : std_logic ;
  signal N_1576 : std_logic ;
  signal N_4660 : std_logic ;
  signal N_1493 : std_logic ;
  signal N_1547 : std_logic ;
  signal N_4661 : std_logic ;
  signal N_1399 : std_logic ;
  signal N_1575 : std_logic ;
  signal N_4662 : std_logic ;
  signal N_1491 : std_logic ;
  signal N_1546 : std_logic ;
  signal N_4663 : std_logic ;
  signal N_1397 : std_logic ;
  signal N_1574 : std_logic ;
  signal N_4664 : std_logic ;
  signal N_1489 : std_logic ;
  signal N_1545 : std_logic ;
  signal N_4665 : std_logic ;
  signal N_1395 : std_logic ;
  signal N_1573 : std_logic ;
  signal N_4666 : std_logic ;
  signal N_1487 : std_logic ;
  signal N_1544 : std_logic ;
  signal N_4667 : std_logic ;
  signal N_1393 : std_logic ;
  signal N_1572 : std_logic ;
  signal N_4668 : std_logic ;
  signal N_1485 : std_logic ;
  signal N_1543 : std_logic ;
  signal N_4669 : std_logic ;
  signal N_1391 : std_logic ;
  signal N_1571 : std_logic ;
  signal N_4670 : std_logic ;
  signal N_1483 : std_logic ;
  signal N_1542 : std_logic ;
  signal N_4671 : std_logic ;
  signal N_1389 : std_logic ;
  signal N_1570 : std_logic ;
  signal N_4672 : std_logic ;
  signal N_1481 : std_logic ;
  signal N_1541 : std_logic ;
  signal N_4673 : std_logic ;
  signal N_1387 : std_logic ;
  signal N_1569 : std_logic ;
  signal N_4674 : std_logic ;
  signal N_1479 : std_logic ;
  signal N_1540 : std_logic ;
  signal N_4675 : std_logic ;
  signal N_1385 : std_logic ;
  signal N_1568 : std_logic ;
  signal N_4676 : std_logic ;
  signal N_1477 : std_logic ;
  signal N_1539 : std_logic ;
  signal N_4677 : std_logic ;
  signal N_1383 : std_logic ;
  signal N_1567 : std_logic ;
  signal N_4678 : std_logic ;
  signal N_1475 : std_logic ;
  signal N_1538 : std_logic ;
  signal N_4679 : std_logic ;
  signal N_1381 : std_logic ;
  signal N_1566 : std_logic ;
  signal N_4680 : std_logic ;
  signal N_1473 : std_logic ;
  signal N_1537 : std_logic ;
  signal N_4681 : std_logic ;
  signal N_1379 : std_logic ;
  signal N_1565 : std_logic ;
  signal N_4682 : std_logic ;
  signal N_1471 : std_logic ;
  signal N_1536 : std_logic ;
  signal N_4683 : std_logic ;
  signal N_1469 : std_logic ;
  signal N_1535 : std_logic ;
  signal N_4684 : std_logic ;
  signal N_1467 : std_logic ;
  signal N_1534 : std_logic ;
  signal N_4685 : std_logic ;
  signal N_1465 : std_logic ;
  signal N_1533 : std_logic ;
  signal N_4686 : std_logic ;
  signal N_1463 : std_logic ;
  signal N_1532 : std_logic ;
  signal N_4687 : std_logic ;
  signal N_1461 : std_logic ;
  signal N_1531 : std_logic ;
  signal N_4688 : std_logic ;
  signal N_1459 : std_logic ;
  signal N_1530 : std_logic ;
  signal N_4689 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_0 : std_logic ;
  signal R1IN_ADD_1_1_AXB_0 : std_logic ;
  signal N_4690 : std_logic ;
  signal N_1457 : std_logic ;
  signal N_1529 : std_logic ;
  signal N_4691 : std_logic ;
  signal N_1455 : std_logic ;
  signal N_1528 : std_logic ;
  signal N_4692 : std_logic ;
  signal N_1453 : std_logic ;
  signal N_1527 : std_logic ;
  signal N_4693 : std_logic ;
  signal N_1451 : std_logic ;
  signal N_1526 : std_logic ;
  signal N_4694 : std_logic ;
  signal N_1449 : std_logic ;
  signal N_1525 : std_logic ;
  signal N_4695 : std_logic ;
  signal N_1447 : std_logic ;
  signal N_1524 : std_logic ;
  signal N_4696 : std_logic ;
  signal N_1445 : std_logic ;
  signal N_1523 : std_logic ;
  signal N_4697 : std_logic ;
  signal N_4698 : std_logic ;
  signal N_4699 : std_logic ;
  signal N_4700 : std_logic ;
  signal N_4701 : std_logic ;
  signal N_4702 : std_logic ;
  signal N_4703 : std_logic ;
  signal N_4704 : std_logic ;
  signal N_4705 : std_logic ;
  signal N_4706 : std_logic ;
  signal N_4707 : std_logic ;
  signal N_4708 : std_logic ;
  signal N_4709 : std_logic ;
  signal N_4710 : std_logic ;
  signal N_4711 : std_logic ;
  signal N_4712 : std_logic ;
  signal N_4713 : std_logic ;
  signal N_4714 : std_logic ;
  signal N_4715 : std_logic ;
  signal N_4716 : std_logic ;
  signal N_4717 : std_logic ;
  signal N_4718 : std_logic ;
  signal N_4719 : std_logic ;
  signal N_4720 : std_logic ;
  signal N_4721 : std_logic ;
  signal N_4722 : std_logic ;
  signal N_4723 : std_logic ;
  signal N_4724 : std_logic ;
  signal N_4725 : std_logic ;
  signal N_4726 : std_logic ;
  signal N_4727 : std_logic ;
  signal N_4728 : std_logic ;
  signal N_4729 : std_logic ;
  signal N_4730 : std_logic ;
  signal N_4731 : std_logic ;
  signal N_4732 : std_logic ;
  signal N_4733 : std_logic ;
  signal N_4734 : std_logic ;
  signal N_4735 : std_logic ;
  signal N_4736 : std_logic ;
  signal N_4737 : std_logic ;
  signal N_4738 : std_logic ;
  signal N_4739 : std_logic ;
  signal N_4740 : std_logic ;
  signal N_4741 : std_logic ;
  signal N_4742 : std_logic ;
  signal N_4743 : std_logic ;
  signal N_4744 : std_logic ;
  signal N_4745 : std_logic ;
  signal N_4746 : std_logic ;
  signal N_4747 : std_logic ;
  signal N_4748 : std_logic ;
  signal N_4749 : std_logic ;
  signal N_4750 : std_logic ;
  signal N_4751 : std_logic ;
  signal N_4752 : std_logic ;
  signal N_4753 : std_logic ;
  signal N_4754 : std_logic ;
  signal N_4755 : std_logic ;
  signal N_4756 : std_logic ;
  signal N_4757 : std_logic ;
  signal N_4758 : std_logic ;
  signal R1IN_3_ADD_1_RETO : std_logic ;
  signal N_4759 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_0 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_0 : std_logic ;
  signal N_4760 : std_logic ;
  signal N_4761 : std_logic ;
  signal N_4762 : std_logic ;
  signal N_4763 : std_logic ;
  signal N_4764 : std_logic ;
  signal N_4765 : std_logic ;
  signal N_4766 : std_logic ;
  signal N_4767 : std_logic ;
  signal N_4768 : std_logic ;
  signal N_4769 : std_logic ;
  signal N_4770 : std_logic ;
  signal N_4771 : std_logic ;
  signal N_4772 : std_logic ;
  signal N_4773 : std_logic ;
  signal N_4774 : std_logic ;
  signal N_4775 : std_logic ;
  signal N_4776 : std_logic ;
  signal N_4777 : std_logic ;
  signal N_4778 : std_logic ;
  signal N_4779 : std_logic ;
  signal N_4780 : std_logic ;
  signal N_4781 : std_logic ;
  signal N_4782 : std_logic ;
  signal N_4783 : std_logic ;
  signal N_4784 : std_logic ;
  signal N_4785 : std_logic ;
  signal N_4786 : std_logic ;
  signal N_4787 : std_logic ;
  signal N_4788 : std_logic ;
  signal N_4789 : std_logic ;
  signal N_4790 : std_logic ;
  signal N_4791 : std_logic ;
  signal N_4792 : std_logic ;
  signal N_4793 : std_logic ;
  signal N_4794 : std_logic ;
  signal N_4795 : std_logic ;
  signal N_4796 : std_logic ;
  signal N_4797 : std_logic ;
  signal N_4798 : std_logic ;
  signal N_4799 : std_logic ;
  signal N_4800 : std_logic ;
  signal N_4801 : std_logic ;
  signal N_4802 : std_logic ;
  signal N_4803 : std_logic ;
  signal N_4804 : std_logic ;
  signal N_4805 : std_logic ;
  signal N_4806 : std_logic ;
  signal N_4807 : std_logic ;
  signal N_4808 : std_logic ;
  signal N_4809 : std_logic ;
  signal N_4810 : std_logic ;
  signal N_4811 : std_logic ;
  signal N_4812 : std_logic ;
  signal N_4813 : std_logic ;
  signal N_4814 : std_logic ;
  signal N_4815 : std_logic ;
  signal N_4816 : std_logic ;
  signal N_4817 : std_logic ;
  signal N_4818 : std_logic ;
  signal N_4819 : std_logic ;
  signal N_4820 : std_logic ;
  signal N_4821 : std_logic ;
  signal N_4822 : std_logic ;
  signal N_4823 : std_logic ;
  signal N_4824 : std_logic ;
  signal N_4825 : std_logic ;
  signal N_4826 : std_logic ;
  signal N_4827 : std_logic ;
  signal N_4828 : std_logic ;
  signal N_4829 : std_logic ;
  signal N_4830 : std_logic ;
  signal R1IN_4_ADD_2_0_RETO : std_logic ;
  signal R1IN_4_4_ADD_2_RETO : std_logic ;
  signal N_4831 : std_logic ;
  signal N_4880 : std_logic ;
  signal N_4881 : std_logic ;
  signal N_4882 : std_logic ;
  signal N_4883 : std_logic ;
  signal N_4884 : std_logic ;
  signal N_4885 : std_logic ;
  signal N_4886 : std_logic ;
  signal N_4887 : std_logic ;
  signal N_4888 : std_logic ;
  signal N_4889 : std_logic ;
  signal N_4890 : std_logic ;
  signal N_4891 : std_logic ;
  signal N_4892 : std_logic ;
  signal N_4893 : std_logic ;
  signal N_4894 : std_logic ;
  signal N_4895 : std_logic ;
  signal N_4896 : std_logic ;
  signal N_4897 : std_logic ;
  signal N_4898 : std_logic ;
  signal N_4899 : std_logic ;
  signal N_4900 : std_logic ;
  signal N_4901 : std_logic ;
  signal N_4902 : std_logic ;
  signal N_4903 : std_logic ;
  signal N_4904 : std_logic ;
  signal N_4905 : std_logic ;
  signal N_4906 : std_logic ;
  signal N_4907 : std_logic ;
  signal N_4908 : std_logic ;
  signal N_4909 : std_logic ;
  signal N_4910 : std_logic ;
  signal N_4911 : std_logic ;
  signal N_4912 : std_logic ;
  signal N_4913 : std_logic ;
  signal N_4914 : std_logic ;
  signal N_4915 : std_logic ;
  signal N_4916 : std_logic ;
  signal N_4917 : std_logic ;
  signal N_4918 : std_logic ;
  signal N_4919 : std_logic ;
  signal N_4920 : std_logic ;
  signal N_4921 : std_logic ;
  signal N_4922 : std_logic ;
  signal N_4923 : std_logic ;
  signal N_4924 : std_logic ;
  signal N_4925 : std_logic ;
  signal N_4926 : std_logic ;
  signal N_4927 : std_logic ;
  signal N_4928 : std_logic ;
  signal N_4929 : std_logic ;
  signal N_4930 : std_logic ;
  signal N_4931 : std_logic ;
  signal N_4932 : std_logic ;
  signal N_4933 : std_logic ;
  signal N_4934 : std_logic ;
  signal N_4935 : std_logic ;
  signal N_4936 : std_logic ;
  signal N_4937 : std_logic ;
  signal N_4938 : std_logic ;
  signal N_4939 : std_logic ;
  signal N_4940 : std_logic ;
  signal N_4941 : std_logic ;
  signal N_4942 : std_logic ;
  signal N_4943 : std_logic ;
  signal N_4944 : std_logic ;
  signal N_4945 : std_logic ;
  signal N_4946 : std_logic ;
  signal N_4947 : std_logic ;
  signal N_4948 : std_logic ;
  signal N_4949 : std_logic ;
  signal N_4950 : std_logic ;
  signal N_4951 : std_logic ;
  signal N_4952 : std_logic ;
  signal N_4953 : std_logic ;
  signal N_4954 : std_logic ;
  signal N_4955 : std_logic ;
  signal N_4956 : std_logic ;
  signal N_4957 : std_logic ;
  signal N_4958 : std_logic ;
  signal N_4959 : std_logic ;
  signal N_4960 : std_logic ;
  signal N_4961 : std_logic ;
  signal N_4962 : std_logic ;
  signal N_4963 : std_logic ;
  signal N_4964 : std_logic ;
  signal N_4965 : std_logic ;
  signal N_4966 : std_logic ;
  signal N_4967 : std_logic ;
  signal N_4968 : std_logic ;
  signal N_4969 : std_logic ;
  signal N_4970 : std_logic ;
  signal N_4971 : std_logic ;
  signal N_4972 : std_logic ;
  signal N_4973 : std_logic ;
  signal N_4974 : std_logic ;
  signal N_4975 : std_logic ;
  signal N_4976 : std_logic ;
  signal N_4977 : std_logic ;
  signal N_4978 : std_logic ;
  signal N_4979 : std_logic ;
  signal N_4980 : std_logic ;
  signal N_4981 : std_logic ;
  signal N_4982 : std_logic ;
  signal N_4983 : std_logic ;
  signal N_4984 : std_logic ;
  signal N_4985 : std_logic ;
  signal N_4986 : std_logic ;
  signal N_4987 : std_logic ;
  signal N_4988 : std_logic ;
  signal N_4989 : std_logic ;
  signal N_4990 : std_logic ;
  signal N_4991 : std_logic ;
  signal N_4992 : std_logic ;
  signal N_4993 : std_logic ;
  signal N_4994 : std_logic ;
  signal N_4995 : std_logic ;
  signal N_4996 : std_logic ;
  signal N_4997 : std_logic ;
  signal N_4998 : std_logic ;
  signal N_4999 : std_logic ;
  signal N_5000 : std_logic ;
  signal N_5001 : std_logic ;
  signal N_5002 : std_logic ;
  signal N_5003 : std_logic ;
  signal N_5004 : std_logic ;
  signal N_5005 : std_logic ;
  signal N_5006 : std_logic ;
  signal N_5007 : std_logic ;
  signal N_5008 : std_logic ;
  signal R1IN_4_ADD_2_1_RETO : std_logic ;
  signal N_5009 : std_logic ;
  signal N_5010 : std_logic ;
  signal N_5011 : std_logic ;
  signal N_5012 : std_logic ;
  signal N_5013 : std_logic ;
  signal N_5014 : std_logic ;
  signal N_5015 : std_logic ;
  signal N_5016 : std_logic ;
  signal N_5017 : std_logic ;
  signal N_5018 : std_logic ;
  signal N_5019 : std_logic ;
  signal N_5020 : std_logic ;
  signal N_5021 : std_logic ;
  signal N_5022 : std_logic ;
  signal N_5023 : std_logic ;
  signal N_5024 : std_logic ;
  signal N_5025 : std_logic ;
  signal N_5026 : std_logic ;
  signal N_5027 : std_logic ;
  signal N_5028 : std_logic ;
  signal N_5029 : std_logic ;
  signal N_5030 : std_logic ;
  signal N_5031 : std_logic ;
  signal N_5032 : std_logic ;
  signal N_5033 : std_logic ;
  signal N_5034 : std_logic ;
  signal N_5035 : std_logic ;
  signal N_5036 : std_logic ;
  signal N_5037 : std_logic ;
  signal N_5038 : std_logic ;
  signal N_5039 : std_logic ;
  signal N_5040 : std_logic ;
  signal N_5041 : std_logic ;
  signal N_5042 : std_logic ;
  signal N_5043 : std_logic ;
  signal N_5044 : std_logic ;
  signal N_5045 : std_logic ;
  signal N_5046 : std_logic ;
  signal N_5047 : std_logic ;
  signal N_5048 : std_logic ;
  signal N_5049 : std_logic ;
  signal N_5050 : std_logic ;
  signal N_5051 : std_logic ;
  signal N_5052 : std_logic ;
  signal N_5053 : std_logic ;
  signal N_5054 : std_logic ;
  signal N_5055 : std_logic ;
  signal N_5056 : std_logic ;
  signal N_5057 : std_logic ;
  signal N_5058 : std_logic ;
  signal N_5059 : std_logic ;
  signal N_5060 : std_logic ;
  signal N_5061 : std_logic ;
  signal N_5062 : std_logic ;
  signal N_5063 : std_logic ;
  signal N_5064 : std_logic ;
  signal N_5065 : std_logic ;
  signal N_5066 : std_logic ;
  signal N_5067 : std_logic ;
  signal N_5068 : std_logic ;
  signal N_5069 : std_logic ;
  signal N_5070 : std_logic ;
  signal N_5071 : std_logic ;
  signal N_5072 : std_logic ;
  signal N_5073 : std_logic ;
  signal N_5074 : std_logic ;
  signal N_5075 : std_logic ;
  signal N_5076 : std_logic ;
  signal N_5077 : std_logic ;
  signal N_5078 : std_logic ;
  signal N_5079 : std_logic ;
  signal N_5080 : std_logic ;
  signal N_5081 : std_logic ;
  signal R1IN_3_ADD_1 : std_logic ;
  signal R1IN_3_ADD_1_RETO_0 : std_logic ;
  signal N_5082 : std_logic ;
  signal N_5083 : std_logic ;
  signal N_5084 : std_logic ;
  signal N_5085 : std_logic ;
  signal N_5086 : std_logic ;
  signal N_5087 : std_logic ;
  signal N_5088 : std_logic ;
  signal N_5089 : std_logic ;
  signal N_5090 : std_logic ;
  signal N_5091 : std_logic ;
  signal N_5092 : std_logic ;
  signal N_5093 : std_logic ;
  signal N_5094 : std_logic ;
  signal N_5095 : std_logic ;
  signal N_5096 : std_logic ;
  signal N_5097 : std_logic ;
  signal N_5098 : std_logic ;
  signal N_5099 : std_logic ;
  signal N_5100 : std_logic ;
  signal N_5101 : std_logic ;
  signal N_5102 : std_logic ;
  signal N_5103 : std_logic ;
  signal N_5104 : std_logic ;
  signal N_5105 : std_logic ;
  signal N_5106 : std_logic ;
  signal N_5107 : std_logic ;
  signal N_5108 : std_logic ;
  signal N_5109 : std_logic ;
  signal N_5110 : std_logic ;
  signal N_5111 : std_logic ;
  signal N_5112 : std_logic ;
  signal N_5113 : std_logic ;
  signal N_5114 : std_logic ;
  signal N_5115 : std_logic ;
  signal N_5116 : std_logic ;
  signal N_5117 : std_logic ;
  signal N_5118 : std_logic ;
  signal N_5119 : std_logic ;
  signal N_5120 : std_logic ;
  signal N_5121 : std_logic ;
  signal N_5122 : std_logic ;
  signal N_5123 : std_logic ;
  signal N_5124 : std_logic ;
  signal N_5125 : std_logic ;
  signal N_5126 : std_logic ;
  signal N_5127 : std_logic ;
  signal N_5128 : std_logic ;
  signal N_5129 : std_logic ;
  signal N_5130 : std_logic ;
  signal N_5131 : std_logic ;
  signal N_5132 : std_logic ;
  signal N_5133 : std_logic ;
  signal N_5134 : std_logic ;
  signal N_5135 : std_logic ;
  signal N_5136 : std_logic ;
  signal N_5137 : std_logic ;
  signal N_5138 : std_logic ;
  signal N_5139 : std_logic ;
  signal N_5140 : std_logic ;
  signal N_5141 : std_logic ;
  signal N_5142 : std_logic ;
  signal N_5143 : std_logic ;
  signal N_5144 : std_logic ;
  signal N_5145 : std_logic ;
  signal N_5146 : std_logic ;
  signal N_5147 : std_logic ;
  signal N_5148 : std_logic ;
  signal N_5149 : std_logic ;
  signal N_5150 : std_logic ;
  signal N_5151 : std_logic ;
  signal N_5152 : std_logic ;
  signal R1IN_4_4_ADD_2 : std_logic ;
  signal R1IN_4_4_ADD_2_RETO_0 : std_logic ;
  signal N_5153 : std_logic ;
  signal R1IN_2_ADD_1_AXB_1 : std_logic ;
  signal R1IN_2_ADD_1_CRY_0 : std_logic ;
  signal R1IN_2_ADD_1_AXB_2 : std_logic ;
  signal R1IN_2_ADD_1_CRY_1 : std_logic ;
  signal R1IN_2_ADD_1_AXB_3 : std_logic ;
  signal R1IN_2_ADD_1_CRY_2 : std_logic ;
  signal R1IN_2_ADD_1_AXB_4 : std_logic ;
  signal R1IN_2_ADD_1_CRY_3 : std_logic ;
  signal R1IN_2_ADD_1_AXB_5 : std_logic ;
  signal R1IN_2_ADD_1_CRY_4 : std_logic ;
  signal R1IN_2_ADD_1_AXB_6 : std_logic ;
  signal R1IN_2_ADD_1_CRY_5 : std_logic ;
  signal R1IN_2_ADD_1_AXB_7 : std_logic ;
  signal R1IN_2_ADD_1_CRY_6 : std_logic ;
  signal R1IN_2_ADD_1_AXB_8 : std_logic ;
  signal R1IN_2_ADD_1_CRY_7 : std_logic ;
  signal R1IN_2_ADD_1_AXB_9 : std_logic ;
  signal R1IN_2_ADD_1_CRY_8 : std_logic ;
  signal R1IN_2_ADD_1_AXB_10 : std_logic ;
  signal R1IN_2_ADD_1_CRY_9 : std_logic ;
  signal R1IN_2_ADD_1_AXB_11 : std_logic ;
  signal R1IN_2_ADD_1_CRY_10 : std_logic ;
  signal R1IN_2_ADD_1_AXB_12 : std_logic ;
  signal R1IN_2_ADD_1_CRY_11 : std_logic ;
  signal R1IN_2_ADD_1_AXB_13 : std_logic ;
  signal R1IN_2_ADD_1_CRY_12 : std_logic ;
  signal R1IN_2_ADD_1_AXB_14 : std_logic ;
  signal R1IN_2_ADD_1_CRY_13 : std_logic ;
  signal R1IN_2_ADD_1_AXB_15 : std_logic ;
  signal R1IN_2_ADD_1_CRY_14 : std_logic ;
  signal R1IN_2_ADD_1_AXB_16 : std_logic ;
  signal R1IN_2_ADD_1_CRY_15 : std_logic ;
  signal R1IN_2_ADD_1_AXB_17 : std_logic ;
  signal R1IN_2_ADD_1_CRY_16 : std_logic ;
  signal R1IN_2_ADD_1_AXB_18 : std_logic ;
  signal R1IN_2_ADD_1_CRY_17 : std_logic ;
  signal R1IN_2_ADD_1_AXB_19 : std_logic ;
  signal R1IN_2_ADD_1_CRY_18 : std_logic ;
  signal R1IN_2_ADD_1_AXB_20 : std_logic ;
  signal R1IN_2_ADD_1_CRY_19 : std_logic ;
  signal R1IN_2_ADD_1_AXB_21 : std_logic ;
  signal R1IN_2_ADD_1_CRY_20 : std_logic ;
  signal R1IN_2_ADD_1_AXB_22 : std_logic ;
  signal R1IN_2_ADD_1_CRY_21 : std_logic ;
  signal R1IN_2_ADD_1_AXB_23 : std_logic ;
  signal R1IN_2_ADD_1_CRY_22 : std_logic ;
  signal R1IN_2_ADD_1_AXB_24 : std_logic ;
  signal R1IN_2_ADD_1_CRY_23 : std_logic ;
  signal R1IN_2_ADD_1_AXB_25 : std_logic ;
  signal R1IN_2_ADD_1_CRY_24 : std_logic ;
  signal R1IN_2_ADD_1_AXB_26 : std_logic ;
  signal R1IN_2_ADD_1_CRY_25 : std_logic ;
  signal R1IN_2_ADD_1_AXB_27 : std_logic ;
  signal R1IN_2_ADD_1_CRY_26 : std_logic ;
  signal R1IN_2_ADD_1_AXB_28 : std_logic ;
  signal R1IN_2_ADD_1_CRY_27 : std_logic ;
  signal R1IN_2_ADD_1_AXB_29 : std_logic ;
  signal R1IN_2_ADD_1_CRY_28 : std_logic ;
  signal R1IN_2_ADD_1_AXB_30 : std_logic ;
  signal R1IN_2_ADD_1_CRY_29 : std_logic ;
  signal R1IN_2_ADD_1_AXB_31 : std_logic ;
  signal R1IN_2_ADD_1_CRY_30 : std_logic ;
  signal R1IN_2_ADD_1_AXB_32 : std_logic ;
  signal R1IN_2_ADD_1_CRY_31 : std_logic ;
  signal R1IN_2_ADD_1_AXB_33 : std_logic ;
  signal R1IN_2_ADD_1_CRY_32 : std_logic ;
  signal R1IN_2_ADD_1_AXB_34 : std_logic ;
  signal R1IN_2_ADD_1_CRY_33 : std_logic ;
  signal R1IN_2_ADD_1_AXB_35 : std_logic ;
  signal R1IN_2_ADD_1_CRY_34 : std_logic ;
  signal R1IN_2_ADD_1_AXB_36 : std_logic ;
  signal R1IN_2_ADD_1_CRY_35 : std_logic ;
  signal R1IN_2_ADD_1_AXB_37 : std_logic ;
  signal R1IN_2_ADD_1_CRY_36 : std_logic ;
  signal R1IN_2_ADD_1_AXB_38 : std_logic ;
  signal R1IN_2_ADD_1_CRY_37 : std_logic ;
  signal R1IN_2_ADD_1_AXB_39 : std_logic ;
  signal R1IN_2_ADD_1_CRY_38 : std_logic ;
  signal R1IN_2_ADD_1_AXB_40 : std_logic ;
  signal R1IN_2_ADD_1_CRY_39 : std_logic ;
  signal R1IN_2_ADD_1_AXB_41 : std_logic ;
  signal R1IN_2_ADD_1_CRY_40 : std_logic ;
  signal R1IN_2_ADD_1_AXB_42 : std_logic ;
  signal R1IN_2_ADD_1_CRY_41 : std_logic ;
  signal R1IN_2_ADD_1_CRY_42 : std_logic ;
  signal R1IN_2_ADD_1_AXB_43 : std_logic ;
  signal N_1 : std_logic ;
  signal N_2 : std_logic ;
  signal N_3 : std_logic ;
  signal N_4 : std_logic ;
  signal N_5 : std_logic ;
  signal N_6 : std_logic ;
  signal N_7 : std_logic ;
  signal N_8 : std_logic ;
  signal N_9 : std_logic ;
  signal N_10 : std_logic ;
  signal N_11 : std_logic ;
  signal N_12 : std_logic ;
  signal N_13 : std_logic ;
  signal N_14 : std_logic ;
  signal N_15 : std_logic ;
  signal N_16 : std_logic ;
  signal N_17 : std_logic ;
  signal N_18 : std_logic ;
  signal N_19 : std_logic ;
  signal N_20 : std_logic ;
  signal N_21 : std_logic ;
  signal N_22 : std_logic ;
  signal N_23 : std_logic ;
  signal N_24 : std_logic ;
  signal N_25 : std_logic ;
  signal N_26 : std_logic ;
  signal N_27 : std_logic ;
  signal N_28 : std_logic ;
  signal N_29 : std_logic ;
  signal N_30 : std_logic ;
  signal N_31 : std_logic ;
  signal N_32 : std_logic ;
  signal N_33 : std_logic ;
  signal N_34 : std_logic ;
  signal N_35 : std_logic ;
  signal N_36 : std_logic ;
  signal N_37 : std_logic ;
  signal N_38 : std_logic ;
  signal N_39 : std_logic ;
  signal N_40 : std_logic ;
  signal N_41 : std_logic ;
  signal N_42 : std_logic ;
  signal N_43 : std_logic ;
  signal N_44 : std_logic ;
  signal N_45 : std_logic ;
  signal N_46 : std_logic ;
  signal N_47 : std_logic ;
  signal N_48 : std_logic ;
  signal N_49 : std_logic ;
  signal N_50 : std_logic ;
  signal N_51 : std_logic ;
  signal N_52 : std_logic ;
  signal N_53 : std_logic ;
  signal N_54 : std_logic ;
  signal N_55 : std_logic ;
  signal N_56 : std_logic ;
  signal N_57 : std_logic ;
  signal N_58 : std_logic ;
  signal N_59 : std_logic ;
  signal N_60 : std_logic ;
  signal N_61 : std_logic ;
  signal N_62 : std_logic ;
  signal N_63 : std_logic ;
  signal N_64 : std_logic ;
  signal N_65 : std_logic ;
  signal N_66 : std_logic ;
  signal N_67 : std_logic ;
  signal N_68 : std_logic ;
  signal N_69 : std_logic ;
  signal N_70 : std_logic ;
  signal N_71 : std_logic ;
  signal N_72 : std_logic ;
  signal R1IN_2_ADD_1_RETO : std_logic ;
  signal N_73 : std_logic ;
  signal R1IN_4_ADD_1_AXB_1 : std_logic ;
  signal R1IN_4_ADD_1_CRY_0 : std_logic ;
  signal R1IN_4_ADD_1_AXB_2 : std_logic ;
  signal R1IN_4_ADD_1_CRY_1 : std_logic ;
  signal R1IN_4_ADD_1_AXB_3 : std_logic ;
  signal R1IN_4_ADD_1_CRY_2 : std_logic ;
  signal R1IN_4_ADD_1_AXB_4 : std_logic ;
  signal R1IN_4_ADD_1_CRY_3 : std_logic ;
  signal R1IN_4_ADD_1_AXB_5 : std_logic ;
  signal R1IN_4_ADD_1_CRY_4 : std_logic ;
  signal R1IN_4_ADD_1_AXB_6 : std_logic ;
  signal R1IN_4_ADD_1_CRY_5 : std_logic ;
  signal R1IN_4_ADD_1_AXB_7 : std_logic ;
  signal R1IN_4_ADD_1_CRY_6 : std_logic ;
  signal R1IN_4_ADD_1_AXB_8 : std_logic ;
  signal R1IN_4_ADD_1_CRY_7 : std_logic ;
  signal R1IN_4_ADD_1_AXB_9 : std_logic ;
  signal R1IN_4_ADD_1_CRY_8 : std_logic ;
  signal R1IN_4_ADD_1_AXB_10 : std_logic ;
  signal R1IN_4_ADD_1_CRY_9 : std_logic ;
  signal R1IN_4_ADD_1_AXB_11 : std_logic ;
  signal R1IN_4_ADD_1_CRY_10 : std_logic ;
  signal R1IN_4_ADD_1_AXB_12 : std_logic ;
  signal R1IN_4_ADD_1_CRY_11 : std_logic ;
  signal R1IN_4_ADD_1_AXB_13 : std_logic ;
  signal R1IN_4_ADD_1_CRY_12 : std_logic ;
  signal R1IN_4_ADD_1_AXB_14 : std_logic ;
  signal R1IN_4_ADD_1_CRY_13 : std_logic ;
  signal R1IN_4_ADD_1_AXB_15 : std_logic ;
  signal R1IN_4_ADD_1_CRY_14 : std_logic ;
  signal R1IN_4_ADD_1_AXB_16 : std_logic ;
  signal R1IN_4_ADD_1_CRY_15 : std_logic ;
  signal R1IN_4_ADD_1_AXB_17 : std_logic ;
  signal R1IN_4_ADD_1_CRY_16 : std_logic ;
  signal R1IN_4_ADD_1_AXB_18 : std_logic ;
  signal R1IN_4_ADD_1_CRY_17 : std_logic ;
  signal R1IN_4_ADD_1_AXB_19 : std_logic ;
  signal R1IN_4_ADD_1_CRY_18 : std_logic ;
  signal R1IN_4_ADD_1_AXB_20 : std_logic ;
  signal R1IN_4_ADD_1_CRY_19 : std_logic ;
  signal R1IN_4_ADD_1_AXB_21 : std_logic ;
  signal R1IN_4_ADD_1_CRY_20 : std_logic ;
  signal R1IN_4_ADD_1_AXB_22 : std_logic ;
  signal R1IN_4_ADD_1_CRY_21 : std_logic ;
  signal R1IN_4_ADD_1_AXB_23 : std_logic ;
  signal R1IN_4_ADD_1_CRY_22 : std_logic ;
  signal R1IN_4_ADD_1_AXB_24 : std_logic ;
  signal R1IN_4_ADD_1_CRY_23 : std_logic ;
  signal R1IN_4_ADD_1_AXB_25 : std_logic ;
  signal R1IN_4_ADD_1_CRY_24 : std_logic ;
  signal R1IN_4_ADD_1_AXB_26 : std_logic ;
  signal R1IN_4_ADD_1_CRY_25 : std_logic ;
  signal R1IN_4_ADD_1_AXB_27 : std_logic ;
  signal R1IN_4_ADD_1_CRY_26 : std_logic ;
  signal R1IN_4_ADD_1_AXB_28 : std_logic ;
  signal R1IN_4_ADD_1_CRY_27 : std_logic ;
  signal R1IN_4_ADD_1_AXB_29 : std_logic ;
  signal R1IN_4_ADD_1_CRY_28 : std_logic ;
  signal R1IN_4_ADD_1_AXB_30 : std_logic ;
  signal R1IN_4_ADD_1_CRY_29 : std_logic ;
  signal R1IN_4_ADD_1_AXB_31 : std_logic ;
  signal R1IN_4_ADD_1_CRY_30 : std_logic ;
  signal R1IN_4_ADD_1_AXB_32 : std_logic ;
  signal R1IN_4_ADD_1_CRY_31 : std_logic ;
  signal R1IN_4_ADD_1_AXB_33 : std_logic ;
  signal R1IN_4_ADD_1_CRY_32 : std_logic ;
  signal R1IN_4_ADD_1_AXB_34 : std_logic ;
  signal R1IN_4_ADD_1_CRY_33 : std_logic ;
  signal R1IN_4_ADD_1_AXB_35 : std_logic ;
  signal R1IN_4_ADD_1_CRY_34 : std_logic ;
  signal R1IN_4_ADD_1_AXB_36 : std_logic ;
  signal R1IN_4_ADD_1_CRY_35 : std_logic ;
  signal R1IN_4_ADD_1_AXB_37 : std_logic ;
  signal R1IN_4_ADD_1_CRY_36 : std_logic ;
  signal R1IN_4_ADD_1_AXB_38 : std_logic ;
  signal R1IN_4_ADD_1_CRY_37 : std_logic ;
  signal R1IN_4_ADD_1_AXB_39 : std_logic ;
  signal R1IN_4_ADD_1_CRY_38 : std_logic ;
  signal R1IN_4_ADD_1_AXB_40 : std_logic ;
  signal R1IN_4_ADD_1_CRY_39 : std_logic ;
  signal R1IN_4_ADD_1_AXB_41 : std_logic ;
  signal R1IN_4_ADD_1_CRY_40 : std_logic ;
  signal R1IN_4_ADD_1_AXB_42 : std_logic ;
  signal R1IN_4_ADD_1_CRY_41 : std_logic ;
  signal R1IN_4_ADD_1_CRY_42 : std_logic ;
  signal R1IN_4_ADD_1_AXB_43 : std_logic ;
  signal N_1_0 : std_logic ;
  signal N_2_0 : std_logic ;
  signal N_3_0 : std_logic ;
  signal N_4_0 : std_logic ;
  signal N_5_0 : std_logic ;
  signal N_6_0 : std_logic ;
  signal N_7_0 : std_logic ;
  signal N_8_0 : std_logic ;
  signal N_9_0 : std_logic ;
  signal N_10_0 : std_logic ;
  signal N_11_0 : std_logic ;
  signal N_12_0 : std_logic ;
  signal N_13_0 : std_logic ;
  signal N_14_0 : std_logic ;
  signal N_15_0 : std_logic ;
  signal N_16_0 : std_logic ;
  signal N_17_0 : std_logic ;
  signal N_18_0 : std_logic ;
  signal N_19_0 : std_logic ;
  signal N_20_0 : std_logic ;
  signal N_21_0 : std_logic ;
  signal N_22_0 : std_logic ;
  signal N_23_0 : std_logic ;
  signal N_24_0 : std_logic ;
  signal N_25_0 : std_logic ;
  signal N_26_0 : std_logic ;
  signal N_27_0 : std_logic ;
  signal N_28_0 : std_logic ;
  signal N_29_0 : std_logic ;
  signal N_30_0 : std_logic ;
  signal N_31_0 : std_logic ;
  signal N_32_0 : std_logic ;
  signal N_33_0 : std_logic ;
  signal N_34_0 : std_logic ;
  signal N_35_0 : std_logic ;
  signal N_36_0 : std_logic ;
  signal N_37_0 : std_logic ;
  signal N_38_0 : std_logic ;
  signal N_39_0 : std_logic ;
  signal N_40_0 : std_logic ;
  signal N_41_0 : std_logic ;
  signal N_42_0 : std_logic ;
  signal N_43_0 : std_logic ;
  signal N_44_0 : std_logic ;
  signal N_45_0 : std_logic ;
  signal N_46_0 : std_logic ;
  signal N_47_0 : std_logic ;
  signal N_48_0 : std_logic ;
  signal N_49_0 : std_logic ;
  signal N_50_0 : std_logic ;
  signal N_51_0 : std_logic ;
  signal N_52_0 : std_logic ;
  signal N_53_0 : std_logic ;
  signal NN_4 : std_logic ;
  signal N_54_0 : std_logic ;
begin
R1IN_4_ADD_2_1_AXB_1_Z4370: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(20),
  I1 => R1IN_4_ADD_1_RETO(37),
  O => R1IN_4_ADD_2_1_AXB_1);
R1IN_4_ADD_2_1_AXB_2_Z4371: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(21),
  I1 => R1IN_4_ADD_1_RETO(38),
  O => R1IN_4_ADD_2_1_AXB_2);
R1IN_4_ADD_2_1_AXB_3_Z4372: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(22),
  I1 => R1IN_4_ADD_1_RETO(39),
  O => R1IN_4_ADD_2_1_AXB_3);
R1IN_4_ADD_2_1_AXB_4_Z4373: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(23),
  I1 => R1IN_4_ADD_1_RETO(40),
  O => R1IN_4_ADD_2_1_AXB_4);
R1IN_4_ADD_2_1_AXB_5_Z4374: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(24),
  I1 => R1IN_4_ADD_1_RETO(41),
  O => R1IN_4_ADD_2_1_AXB_5);
R1IN_4_ADD_2_1_AXB_6_Z4375: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(25),
  I1 => R1IN_4_ADD_1_RETO(42),
  O => R1IN_4_ADD_2_1_AXB_6);
R1IN_4_ADD_2_1_AXB_7_Z4376: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(26),
  I1 => R1IN_4_ADD_1_RETO(43),
  O => R1IN_4_ADD_2_1_AXB_7);
R1IN_4_ADD_2_1_AXB_8_Z4377: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(27),
  I1 => R1IN_4_ADD_1_RETO(44),
  O => R1IN_4_ADD_2_1_AXB_8);
R1IN_4_ADD_2_1_AXB_9_Z4378: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(28),
  O => R1IN_4_ADD_2_1_AXB_9);
R1IN_4_ADD_2_1_AXB_10_Z4379: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(29),
  O => R1IN_4_ADD_2_1_AXB_10);
R1IN_4_ADD_2_1_AXB_11_Z4380: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(30),
  O => R1IN_4_ADD_2_1_AXB_11);
R1IN_4_ADD_2_1_AXB_12_Z4381: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(31),
  O => R1IN_4_ADD_2_1_AXB_12);
R1IN_4_ADD_2_1_AXB_13_Z4382: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(32),
  O => R1IN_4_ADD_2_1_AXB_13);
R1IN_4_ADD_2_1_AXB_14_Z4383: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(33),
  O => R1IN_4_ADD_2_1_AXB_14);
R1IN_4_ADD_2_1_AXB_15_Z4384: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(34),
  O => R1IN_4_ADD_2_1_AXB_15);
R1IN_4_ADD_2_1_AXB_16_Z4385: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(35),
  O => R1IN_4_ADD_2_1_AXB_16);
R1IN_4_ADD_2_1_AXB_17_Z4386: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(36),
  O => R1IN_4_ADD_2_1_AXB_17);
R1IN_4_ADD_2_1_AXB_18_Z4387: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(37),
  O => R1IN_4_ADD_2_1_AXB_18);
R1IN_4_ADD_2_1_AXB_19_Z4388: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(38),
  O => R1IN_4_ADD_2_1_AXB_19);
R1IN_4_ADD_2_1_AXB_20_Z4389: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(39),
  O => R1IN_4_ADD_2_1_AXB_20);
R1IN_4_ADD_2_1_AXB_21_Z4390: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(40),
  O => R1IN_4_ADD_2_1_AXB_21);
R1IN_4_ADD_2_1_AXB_22_Z4391: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(41),
  O => R1IN_4_ADD_2_1_AXB_22);
R1IN_4_ADD_2_1_AXB_23_Z4392: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(42),
  O => R1IN_4_ADD_2_1_AXB_23);
R1IN_4_ADD_2_1_AXB_24_Z4393: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(43),
  O => R1IN_4_ADD_2_1_AXB_24);
R1IN_4_ADD_2_1_AXB_25_Z4394: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(44),
  O => R1IN_4_ADD_2_1_AXB_25);
R1IN_4_ADD_2_1_AXB_26_Z4395: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(45),
  O => R1IN_4_ADD_2_1_AXB_26);
R1IN_4_ADD_2_1_AXB_27_Z4396: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(46),
  O => R1IN_4_ADD_2_1_AXB_27);
R1IN_4_ADD_2_1_AXB_28_Z4397: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(47),
  O => R1IN_4_ADD_2_1_AXB_28);
R1IN_4_ADD_2_1_AXB_29_Z4398: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(48),
  O => R1IN_4_ADD_2_1_AXB_29);
R1IN_4_ADD_2_1_AXB_30_Z4399: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(49),
  O => R1IN_4_ADD_2_1_AXB_30);
R1IN_4_ADD_2_1_AXB_31_Z4400: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(50),
  O => R1IN_4_ADD_2_1_AXB_31);
R1IN_4_ADD_2_1_AXB_32_Z4401: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(51),
  O => R1IN_4_ADD_2_1_AXB_32);
R1IN_4_ADD_2_1_AXB_33_Z4402: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(52),
  O => R1IN_4_ADD_2_1_AXB_33);
R1IN_4_ADD_2_1_0_AXB_1_Z4403: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(20),
  I1 => R1IN_4_ADD_1_RETO(37),
  O => R1IN_4_ADD_2_1_0_AXB_1);
R1IN_4_ADD_2_1_0_AXB_2_Z4404: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(21),
  I1 => R1IN_4_ADD_1_RETO(38),
  O => R1IN_4_ADD_2_1_0_AXB_2);
R1IN_4_ADD_2_1_0_AXB_3_Z4405: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(22),
  I1 => R1IN_4_ADD_1_RETO(39),
  O => R1IN_4_ADD_2_1_0_AXB_3);
R1IN_4_ADD_2_1_0_AXB_4_Z4406: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(23),
  I1 => R1IN_4_ADD_1_RETO(40),
  O => R1IN_4_ADD_2_1_0_AXB_4);
R1IN_4_ADD_2_1_0_AXB_5_Z4407: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(24),
  I1 => R1IN_4_ADD_1_RETO(41),
  O => R1IN_4_ADD_2_1_0_AXB_5);
R1IN_4_ADD_2_1_0_AXB_6_Z4408: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(25),
  I1 => R1IN_4_ADD_1_RETO(42),
  O => R1IN_4_ADD_2_1_0_AXB_6);
R1IN_4_ADD_2_1_0_AXB_7_Z4409: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(26),
  I1 => R1IN_4_ADD_1_RETO(43),
  O => R1IN_4_ADD_2_1_0_AXB_7);
R1IN_4_ADD_2_1_0_AXB_8_Z4410: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(27),
  I1 => R1IN_4_ADD_1_RETO(44),
  O => R1IN_4_ADD_2_1_0_AXB_8);
R1IN_4_ADD_2_1_0_AXB_9_Z4411: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(28),
  O => R1IN_4_ADD_2_1_0_AXB_9);
R1IN_4_ADD_2_1_0_AXB_10_Z4412: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(29),
  O => R1IN_4_ADD_2_1_0_AXB_10);
R1IN_4_ADD_2_1_0_AXB_11_Z4413: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(30),
  O => R1IN_4_ADD_2_1_0_AXB_11);
R1IN_4_ADD_2_1_0_AXB_12_Z4414: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(31),
  O => R1IN_4_ADD_2_1_0_AXB_12);
R1IN_4_ADD_2_1_0_AXB_13_Z4415: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(32),
  O => R1IN_4_ADD_2_1_0_AXB_13);
R1IN_4_ADD_2_1_0_AXB_14_Z4416: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(33),
  O => R1IN_4_ADD_2_1_0_AXB_14);
R1IN_4_ADD_2_1_0_AXB_15_Z4417: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(34),
  O => R1IN_4_ADD_2_1_0_AXB_15);
R1IN_4_ADD_2_1_0_AXB_16_Z4418: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(35),
  O => R1IN_4_ADD_2_1_0_AXB_16);
R1IN_4_ADD_2_1_0_AXB_17_Z4419: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(36),
  O => R1IN_4_ADD_2_1_0_AXB_17);
R1IN_4_ADD_2_1_0_AXB_18_Z4420: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(37),
  O => R1IN_4_ADD_2_1_0_AXB_18);
R1IN_4_ADD_2_1_0_AXB_19_Z4421: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(38),
  O => R1IN_4_ADD_2_1_0_AXB_19);
R1IN_4_ADD_2_1_0_AXB_20_Z4422: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(39),
  O => R1IN_4_ADD_2_1_0_AXB_20);
R1IN_4_ADD_2_1_0_AXB_21_Z4423: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(40),
  O => R1IN_4_ADD_2_1_0_AXB_21);
R1IN_4_ADD_2_1_0_AXB_22_Z4424: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(41),
  O => R1IN_4_ADD_2_1_0_AXB_22);
R1IN_4_ADD_2_1_0_AXB_23_Z4425: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(42),
  O => R1IN_4_ADD_2_1_0_AXB_23);
R1IN_4_ADD_2_1_0_AXB_24_Z4426: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(43),
  O => R1IN_4_ADD_2_1_0_AXB_24);
R1IN_4_ADD_2_1_0_AXB_25_Z4427: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(44),
  O => R1IN_4_ADD_2_1_0_AXB_25);
R1IN_4_ADD_2_1_0_AXB_26_Z4428: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(45),
  O => R1IN_4_ADD_2_1_0_AXB_26);
R1IN_4_ADD_2_1_0_AXB_27_Z4429: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(46),
  O => R1IN_4_ADD_2_1_0_AXB_27);
R1IN_4_ADD_2_1_0_AXB_28_Z4430: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(47),
  O => R1IN_4_ADD_2_1_0_AXB_28);
R1IN_4_ADD_2_1_0_AXB_29_Z4431: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(48),
  O => R1IN_4_ADD_2_1_0_AXB_29);
R1IN_4_ADD_2_1_0_AXB_30_Z4432: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(49),
  O => R1IN_4_ADD_2_1_0_AXB_30);
R1IN_4_ADD_2_1_0_AXB_31_Z4433: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(50),
  O => R1IN_4_ADD_2_1_0_AXB_31);
R1IN_4_ADD_2_1_0_AXB_32_Z4434: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(51),
  O => R1IN_4_ADD_2_1_0_AXB_32);
R1IN_4_ADD_2_1_0_AXB_33_Z4435: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(52),
  O => R1IN_4_ADD_2_1_0_AXB_33);
R1IN_ADD_1_1_AXB_1_Z4436: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(33),
  I1 => R1IN_3(33),
  O => R1IN_ADD_1_1_AXB_1);
R1IN_ADD_1_1_AXB_2_Z4437: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(34),
  I1 => R1IN_3(34),
  O => R1IN_ADD_1_1_AXB_2);
R1IN_ADD_1_1_AXB_3_Z4438: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(35),
  I1 => R1IN_3(35),
  O => R1IN_ADD_1_1_AXB_3);
R1IN_ADD_1_1_AXB_4_Z4439: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(36),
  I1 => R1IN_3(36),
  O => R1IN_ADD_1_1_AXB_4);
R1IN_ADD_1_1_AXB_5_Z4440: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(37),
  I1 => R1IN_3(37),
  O => R1IN_ADD_1_1_AXB_5);
R1IN_ADD_1_1_AXB_6_Z4441: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(38),
  I1 => R1IN_3(38),
  O => R1IN_ADD_1_1_AXB_6);
R1IN_ADD_1_1_AXB_7_Z4442: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(39),
  I1 => R1IN_3(39),
  O => R1IN_ADD_1_1_AXB_7);
R1IN_ADD_1_1_AXB_8_Z4443: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(40),
  I1 => R1IN_3(40),
  O => R1IN_ADD_1_1_AXB_8);
R1IN_ADD_1_1_AXB_9_Z4444: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(41),
  I1 => R1IN_3(41),
  O => R1IN_ADD_1_1_AXB_9);
R1IN_ADD_1_1_AXB_10_Z4445: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(42),
  I1 => R1IN_3(42),
  O => R1IN_ADD_1_1_AXB_10);
R1IN_ADD_1_1_AXB_11_Z4446: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(43),
  I1 => R1IN_3(43),
  O => R1IN_ADD_1_1_AXB_11);
R1IN_ADD_1_1_AXB_12_Z4447: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(44),
  I1 => R1IN_3(44),
  O => R1IN_ADD_1_1_AXB_12);
R1IN_ADD_1_1_AXB_13_Z4448: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(45),
  I1 => R1IN_3(45),
  O => R1IN_ADD_1_1_AXB_13);
R1IN_ADD_1_1_AXB_14_Z4449: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(46),
  I1 => R1IN_3(46),
  O => R1IN_ADD_1_1_AXB_14);
R1IN_ADD_1_1_AXB_15_Z4450: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(47),
  I1 => R1IN_3(47),
  O => R1IN_ADD_1_1_AXB_15);
R1IN_ADD_1_1_AXB_16_Z4451: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(48),
  I1 => R1IN_3(48),
  O => R1IN_ADD_1_1_AXB_16);
R1IN_ADD_1_1_AXB_17_Z4452: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(49),
  I1 => R1IN_3(49),
  O => R1IN_ADD_1_1_AXB_17);
R1IN_ADD_1_1_AXB_18_Z4453: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(50),
  I1 => R1IN_3(50),
  O => R1IN_ADD_1_1_AXB_18);
R1IN_ADD_1_1_AXB_19_Z4454: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(51),
  I1 => R1IN_3(51),
  O => R1IN_ADD_1_1_AXB_19);
R1IN_ADD_1_1_AXB_20_Z4455: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(52),
  I1 => R1IN_3(52),
  O => R1IN_ADD_1_1_AXB_20);
R1IN_ADD_1_1_AXB_21_Z4456: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(53),
  I1 => R1IN_3(53),
  O => R1IN_ADD_1_1_AXB_21);
R1IN_ADD_1_1_AXB_22_Z4457: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(54),
  I1 => R1IN_3(54),
  O => R1IN_ADD_1_1_AXB_22);
R1IN_ADD_1_1_AXB_23_Z4458: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(55),
  I1 => R1IN_3(55),
  O => R1IN_ADD_1_1_AXB_23);
R1IN_ADD_1_1_AXB_24_Z4459: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(56),
  I1 => R1IN_3(56),
  O => R1IN_ADD_1_1_AXB_24);
R1IN_ADD_1_1_AXB_25_Z4460: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(57),
  I1 => R1IN_3(57),
  O => R1IN_ADD_1_1_AXB_25);
R1IN_ADD_1_1_AXB_26_Z4461: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(58),
  I1 => R1IN_3(58),
  O => R1IN_ADD_1_1_AXB_26);
R1IN_ADD_1_1_AXB_27_Z4462: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(59),
  I1 => R1IN_3(59),
  O => R1IN_ADD_1_1_AXB_27);
R1IN_ADD_1_1_0_AXB_1_Z4463: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(33),
  I1 => R1IN_3(33),
  O => R1IN_ADD_1_1_0_AXB_1);
R1IN_ADD_1_1_0_AXB_2_Z4464: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(34),
  I1 => R1IN_3(34),
  O => R1IN_ADD_1_1_0_AXB_2);
R1IN_ADD_1_1_0_AXB_3_Z4465: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(35),
  I1 => R1IN_3(35),
  O => R1IN_ADD_1_1_0_AXB_3);
R1IN_ADD_1_1_0_AXB_4_Z4466: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(36),
  I1 => R1IN_3(36),
  O => R1IN_ADD_1_1_0_AXB_4);
R1IN_ADD_1_1_0_AXB_5_Z4467: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(37),
  I1 => R1IN_3(37),
  O => R1IN_ADD_1_1_0_AXB_5);
R1IN_ADD_1_1_0_AXB_6_Z4468: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(38),
  I1 => R1IN_3(38),
  O => R1IN_ADD_1_1_0_AXB_6);
R1IN_ADD_1_1_0_AXB_7_Z4469: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(39),
  I1 => R1IN_3(39),
  O => R1IN_ADD_1_1_0_AXB_7);
R1IN_ADD_1_1_0_AXB_8_Z4470: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(40),
  I1 => R1IN_3(40),
  O => R1IN_ADD_1_1_0_AXB_8);
R1IN_ADD_1_1_0_AXB_9_Z4471: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(41),
  I1 => R1IN_3(41),
  O => R1IN_ADD_1_1_0_AXB_9);
R1IN_ADD_1_1_0_AXB_10_Z4472: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(42),
  I1 => R1IN_3(42),
  O => R1IN_ADD_1_1_0_AXB_10);
R1IN_ADD_1_1_0_AXB_11_Z4473: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(43),
  I1 => R1IN_3(43),
  O => R1IN_ADD_1_1_0_AXB_11);
R1IN_ADD_1_1_0_AXB_12_Z4474: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(44),
  I1 => R1IN_3(44),
  O => R1IN_ADD_1_1_0_AXB_12);
R1IN_ADD_1_1_0_AXB_13_Z4475: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(45),
  I1 => R1IN_3(45),
  O => R1IN_ADD_1_1_0_AXB_13);
R1IN_ADD_1_1_0_AXB_14_Z4476: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(46),
  I1 => R1IN_3(46),
  O => R1IN_ADD_1_1_0_AXB_14);
R1IN_ADD_1_1_0_AXB_15_Z4477: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(47),
  I1 => R1IN_3(47),
  O => R1IN_ADD_1_1_0_AXB_15);
R1IN_ADD_1_1_0_AXB_16_Z4478: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(48),
  I1 => R1IN_3(48),
  O => R1IN_ADD_1_1_0_AXB_16);
R1IN_ADD_1_1_0_AXB_17_Z4479: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(49),
  I1 => R1IN_3(49),
  O => R1IN_ADD_1_1_0_AXB_17);
R1IN_ADD_1_1_0_AXB_18_Z4480: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(50),
  I1 => R1IN_3(50),
  O => R1IN_ADD_1_1_0_AXB_18);
R1IN_ADD_1_1_0_AXB_19_Z4481: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(51),
  I1 => R1IN_3(51),
  O => R1IN_ADD_1_1_0_AXB_19);
R1IN_ADD_1_1_0_AXB_20_Z4482: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(52),
  I1 => R1IN_3(52),
  O => R1IN_ADD_1_1_0_AXB_20);
R1IN_ADD_1_1_0_AXB_21_Z4483: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(53),
  I1 => R1IN_3(53),
  O => R1IN_ADD_1_1_0_AXB_21);
R1IN_ADD_1_1_0_AXB_22_Z4484: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(54),
  I1 => R1IN_3(54),
  O => R1IN_ADD_1_1_0_AXB_22);
R1IN_ADD_1_1_0_AXB_23_Z4485: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(55),
  I1 => R1IN_3(55),
  O => R1IN_ADD_1_1_0_AXB_23);
R1IN_ADD_1_1_0_AXB_24_Z4486: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(56),
  I1 => R1IN_3(56),
  O => R1IN_ADD_1_1_0_AXB_24);
R1IN_ADD_1_1_0_AXB_25_Z4487: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(57),
  I1 => R1IN_3(57),
  O => R1IN_ADD_1_1_0_AXB_25);
R1IN_ADD_1_1_0_AXB_26_Z4488: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(58),
  I1 => R1IN_3(58),
  O => R1IN_ADD_1_1_0_AXB_26);
R1IN_ADD_1_1_0_AXB_27_Z4489: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(59),
  I1 => R1IN_3(59),
  O => R1IN_ADD_1_1_0_AXB_27);
R1IN_ADD_1_1_0_AXB_28_Z4490: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(60),
  I1 => R1IN_3(60),
  O => R1IN_ADD_1_1_0_AXB_28);
R1IN_3_ADD_1_AXB_1_Z4491: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F_RETO(18),
  I1 => R1IN_3_2F_RETO(1),
  O => R1IN_3_ADD_1_AXB_1);
R1IN_3_ADD_1_AXB_2_Z4492: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F_RETO(19),
  I1 => R1IN_3_2F_RETO(2),
  O => R1IN_3_ADD_1_AXB_2);
R1IN_3_ADD_1_AXB_3_Z4493: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F_RETO(20),
  I1 => R1IN_3_2F_RETO(3),
  O => R1IN_3_ADD_1_AXB_3);
R1IN_3_ADD_1_AXB_4_Z4494: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F_RETO(21),
  I1 => R1IN_3_2F_RETO(4),
  O => R1IN_3_ADD_1_AXB_4);
R1IN_3_ADD_1_AXB_5_Z4495: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F_RETO(22),
  I1 => R1IN_3_2F_RETO(5),
  O => R1IN_3_ADD_1_AXB_5);
R1IN_3_ADD_1_AXB_6_Z4496: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F_RETO(23),
  I1 => R1IN_3_2F_RETO(6),
  O => R1IN_3_ADD_1_AXB_6);
R1IN_3_ADD_1_AXB_7_Z4497: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F_RETO(24),
  I1 => R1IN_3_2F_RETO(7),
  O => R1IN_3_ADD_1_AXB_7);
R1IN_3_ADD_1_AXB_8_Z4498: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F_RETO(25),
  I1 => R1IN_3_2F_RETO(8),
  O => R1IN_3_ADD_1_AXB_8);
R1IN_3_ADD_1_AXB_9_Z4499: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F_RETO(26),
  I1 => R1IN_3_2F_RETO(9),
  O => R1IN_3_ADD_1_AXB_9);
R1IN_3_ADD_1_AXB_10_Z4500: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F_RETO(27),
  I1 => R1IN_3_2F_RETO(10),
  O => R1IN_3_ADD_1_AXB_10);
R1IN_3_ADD_1_AXB_11_Z4501: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F_RETO(28),
  I1 => R1IN_3_2F_RETO(11),
  O => R1IN_3_ADD_1_AXB_11);
R1IN_3_ADD_1_AXB_12_Z4502: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F_RETO(29),
  I1 => R1IN_3_2F_RETO(12),
  O => R1IN_3_ADD_1_AXB_12);
R1IN_3_ADD_1_AXB_13_Z4503: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F_RETO(30),
  I1 => R1IN_3_2F_RETO(13),
  O => R1IN_3_ADD_1_AXB_13);
R1IN_3_ADD_1_AXB_14_Z4504: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F_RETO(31),
  I1 => R1IN_3_2F_RETO(14),
  O => R1IN_3_ADD_1_AXB_14);
R1IN_3_ADD_1_AXB_15_Z4505: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F_RETO(32),
  I1 => R1IN_3_2F_RETO(15),
  O => R1IN_3_ADD_1_AXB_15);
R1IN_3_ADD_1_AXB_16_Z4506: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F_RETO(33),
  I1 => R1IN_3_2F_RETO(16),
  O => R1IN_3_ADD_1_AXB_16);
R1IN_3_ADD_1_AXB_17_Z4507: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(17),
  O => R1IN_3_ADD_1_AXB_17);
R1IN_3_ADD_1_AXB_18_Z4508: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(18),
  O => R1IN_3_ADD_1_AXB_18);
R1IN_3_ADD_1_AXB_19_Z4509: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(19),
  O => R1IN_3_ADD_1_AXB_19);
R1IN_3_ADD_1_AXB_20_Z4510: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(20),
  O => R1IN_3_ADD_1_AXB_20);
R1IN_3_ADD_1_AXB_21_Z4511: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(21),
  O => R1IN_3_ADD_1_AXB_21);
R1IN_3_ADD_1_AXB_22_Z4512: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(22),
  O => R1IN_3_ADD_1_AXB_22);
R1IN_3_ADD_1_AXB_23_Z4513: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(23),
  O => R1IN_3_ADD_1_AXB_23);
R1IN_3_ADD_1_AXB_24_Z4514: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(24),
  O => R1IN_3_ADD_1_AXB_24);
R1IN_3_ADD_1_AXB_25_Z4515: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(25),
  O => R1IN_3_ADD_1_AXB_25);
R1IN_3_ADD_1_AXB_26_Z4516: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(26),
  O => R1IN_3_ADD_1_AXB_26);
R1IN_3_ADD_1_AXB_27_Z4517: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(27),
  O => R1IN_3_ADD_1_AXB_27);
R1IN_3_ADD_1_AXB_28_Z4518: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(28),
  O => R1IN_3_ADD_1_AXB_28);
R1IN_3_ADD_1_AXB_29_Z4519: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(29),
  O => R1IN_3_ADD_1_AXB_29);
R1IN_3_ADD_1_AXB_30_Z4520: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(30),
  O => R1IN_3_ADD_1_AXB_30);
R1IN_3_ADD_1_AXB_31_Z4521: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(31),
  O => R1IN_3_ADD_1_AXB_31);
R1IN_3_ADD_1_AXB_32_Z4522: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(32),
  O => R1IN_3_ADD_1_AXB_32);
R1IN_3_ADD_1_AXB_33_Z4523: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(33),
  O => R1IN_3_ADD_1_AXB_33);
R1IN_3_ADD_1_AXB_34_Z4524: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(34),
  O => R1IN_3_ADD_1_AXB_34);
R1IN_3_ADD_1_AXB_35_Z4525: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(35),
  O => R1IN_3_ADD_1_AXB_35);
R1IN_3_ADD_1_AXB_36_Z4526: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(36),
  O => R1IN_3_ADD_1_AXB_36);
R1IN_3_ADD_1_AXB_37_Z4527: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(37),
  O => R1IN_3_ADD_1_AXB_37);
R1IN_3_ADD_1_AXB_38_Z4528: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(38),
  O => R1IN_3_ADD_1_AXB_38);
R1IN_3_ADD_1_AXB_39_Z4529: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(39),
  O => R1IN_3_ADD_1_AXB_39);
R1IN_3_ADD_1_AXB_40_Z4530: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(40),
  O => R1IN_3_ADD_1_AXB_40);
R1IN_3_ADD_1_AXB_41_Z4531: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(41),
  O => R1IN_3_ADD_1_AXB_41);
R1IN_3_ADD_1_AXB_42_Z4532: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(42),
  O => R1IN_3_ADD_1_AXB_42);
R1IN_4_4_ADD_2_AXB_0: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_ADD_1F_RETO_0(0),
  I1 => R1IN_4_4_ADD_2_RETO_0,
  O => R1IN_4_4(17));
R1IN_4_4_ADD_2_AXB_1_Z4534: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F_RETO(18),
  I1 => R1IN_4_4_ADD_1F_RETO(1),
  O => R1IN_4_4_ADD_2_AXB_1);
R1IN_4_4_ADD_2_AXB_2_Z4535: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F_RETO(19),
  I1 => R1IN_4_4_ADD_1F_RETO(2),
  O => R1IN_4_4_ADD_2_AXB_2);
R1IN_4_4_ADD_2_AXB_3_Z4536: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F_RETO(20),
  I1 => R1IN_4_4_ADD_1F_RETO(3),
  O => R1IN_4_4_ADD_2_AXB_3);
R1IN_4_4_ADD_2_AXB_4_Z4537: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F_RETO(21),
  I1 => R1IN_4_4_ADD_1F_RETO(4),
  O => R1IN_4_4_ADD_2_AXB_4);
R1IN_4_4_ADD_2_AXB_5_Z4538: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F_RETO(22),
  I1 => R1IN_4_4_ADD_1F_RETO(5),
  O => R1IN_4_4_ADD_2_AXB_5);
R1IN_4_4_ADD_2_AXB_6_Z4539: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F_RETO(23),
  I1 => R1IN_4_4_ADD_1F_RETO(6),
  O => R1IN_4_4_ADD_2_AXB_6);
R1IN_4_4_ADD_2_AXB_7_Z4540: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F_RETO(24),
  I1 => R1IN_4_4_ADD_1F_RETO(7),
  O => R1IN_4_4_ADD_2_AXB_7);
R1IN_4_4_ADD_2_AXB_8_Z4541: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F_RETO(25),
  I1 => R1IN_4_4_ADD_1F_RETO(8),
  O => R1IN_4_4_ADD_2_AXB_8);
R1IN_4_4_ADD_2_AXB_9_Z4542: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F_RETO(26),
  I1 => R1IN_4_4_ADD_1F_RETO(9),
  O => R1IN_4_4_ADD_2_AXB_9);
R1IN_4_4_ADD_2_AXB_10_Z4543: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F_RETO(27),
  I1 => R1IN_4_4_ADD_1F_RETO(10),
  O => R1IN_4_4_ADD_2_AXB_10);
R1IN_4_4_ADD_2_AXB_11_Z4544: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F_RETO(28),
  I1 => R1IN_4_4_ADD_1F_RETO(11),
  O => R1IN_4_4_ADD_2_AXB_11);
R1IN_4_4_ADD_2_AXB_12_Z4545: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F_RETO(29),
  I1 => R1IN_4_4_ADD_1F_RETO(12),
  O => R1IN_4_4_ADD_2_AXB_12);
R1IN_4_4_ADD_2_AXB_13_Z4546: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F_RETO(30),
  I1 => R1IN_4_4_ADD_1F_RETO(13),
  O => R1IN_4_4_ADD_2_AXB_13);
R1IN_4_4_ADD_2_AXB_14_Z4547: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F_RETO(31),
  I1 => R1IN_4_4_ADD_1F_RETO(14),
  O => R1IN_4_4_ADD_2_AXB_14);
R1IN_4_4_ADD_2_AXB_15_Z4548: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F_RETO(32),
  I1 => R1IN_4_4_ADD_1F_RETO(15),
  O => R1IN_4_4_ADD_2_AXB_15);
R1IN_4_4_ADD_2_AXB_16_Z4549: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F_RETO(33),
  I1 => R1IN_4_4_ADD_1F_RETO(16),
  O => R1IN_4_4_ADD_2_AXB_16);
R1IN_4_4_ADD_2_AXB_17_Z4550: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_4F_RETO(0),
  I1 => R1IN_4_4_ADD_1F_RETO(17),
  O => R1IN_4_4_ADD_2_AXB_17);
R1IN_4_4_ADD_2_AXB_18_Z4551: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_4F_RETO(1),
  I1 => R1IN_4_4_ADD_1F_RETO(18),
  O => R1IN_4_4_ADD_2_AXB_18);
R1IN_4_4_ADD_2_AXB_19_Z4552: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_4F_RETO(2),
  I1 => R1IN_4_4_ADD_1F_RETO(19),
  O => R1IN_4_4_ADD_2_AXB_19);
R1IN_4_4_ADD_2_AXB_20_Z4553: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_4F_RETO(3),
  I1 => R1IN_4_4_ADD_1F_RETO(20),
  O => R1IN_4_4_ADD_2_AXB_20);
R1IN_4_4_ADD_2_AXB_21_Z4554: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_4F_RETO(4),
  I1 => R1IN_4_4_ADD_1F_RETO(21),
  O => R1IN_4_4_ADD_2_AXB_21);
R1IN_4_4_ADD_2_AXB_22_Z4555: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_4F_RETO(5),
  I1 => R1IN_4_4_ADD_1F_RETO(22),
  O => R1IN_4_4_ADD_2_AXB_22);
R1IN_4_4_ADD_2_AXB_23_Z4556: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_4F_RETO(6),
  I1 => R1IN_4_4_ADD_1F_RETO(23),
  O => R1IN_4_4_ADD_2_AXB_23);
R1IN_4_4_ADD_2_AXB_24_Z4557: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_4F_RETO(7),
  I1 => R1IN_4_4_ADD_1F_RETO(24),
  O => R1IN_4_4_ADD_2_AXB_24);
R1IN_4_4_ADD_2_AXB_25_Z4558: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_4F_RETO(8),
  I1 => R1IN_4_4_ADD_1F_RETO(25),
  O => R1IN_4_4_ADD_2_AXB_25);
R1IN_4_4_ADD_2_AXB_26_Z4559: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_4F_RETO(9),
  I1 => R1IN_4_4_ADD_1F_RETO(26),
  O => R1IN_4_4_ADD_2_AXB_26);
R1IN_4_4_ADD_2_AXB_27_Z4560: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_4F_RETO(10),
  I1 => R1IN_4_4_ADD_1F_RETO(27),
  O => R1IN_4_4_ADD_2_AXB_27);
R1IN_4_4_ADD_2_AXB_28_Z4561: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4_4F_RETO(11),
  O => R1IN_4_4_ADD_2_AXB_28);
R1IN_4_4_ADD_2_AXB_29_Z4562: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4_4F_RETO(12),
  O => R1IN_4_4_ADD_2_AXB_29);
R1IN_4_4_ADD_2_AXB_30_Z4563: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4_4F_RETO(13),
  O => R1IN_4_4_ADD_2_AXB_30);
R1IN_4_4_ADD_2_AXB_31_Z4564: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4_4F_RETO(14),
  O => R1IN_4_4_ADD_2_AXB_31);
R1IN_4_4_ADD_2_AXB_32_Z4565: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4_4F_RETO(15),
  O => R1IN_4_4_ADD_2_AXB_32);
R1IN_4_4_ADD_2_AXB_33_Z4566: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4_4F_RETO(16),
  O => R1IN_4_4_ADD_2_AXB_33);
R1IN_4_4_ADD_2_AXB_34_Z4567: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4_4F_RETO(17),
  O => R1IN_4_4_ADD_2_AXB_34);
R1IN_4_4_ADD_2_AXB_35_Z4568: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4_4F_RETO(18),
  O => R1IN_4_4_ADD_2_AXB_35);
R1IN_ADD_2_AXB_1_Z4569: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(18),
  I1 => R1IN_ADD_1(1),
  O => R1IN_ADD_2_AXB_1);
R1IN_ADD_2_AXB_2_Z4570: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(19),
  I1 => R1IN_ADD_1(2),
  O => R1IN_ADD_2_AXB_2);
R1IN_ADD_2_AXB_3_Z4571: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(20),
  I1 => R1IN_ADD_1(3),
  O => R1IN_ADD_2_AXB_3);
R1IN_ADD_2_AXB_4_Z4572: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(21),
  I1 => R1IN_ADD_1(4),
  O => R1IN_ADD_2_AXB_4);
R1IN_ADD_2_AXB_5_Z4573: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(22),
  I1 => R1IN_ADD_1(5),
  O => R1IN_ADD_2_AXB_5);
R1IN_ADD_2_AXB_6_Z4574: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(23),
  I1 => R1IN_ADD_1(6),
  O => R1IN_ADD_2_AXB_6);
R1IN_ADD_2_AXB_7_Z4575: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(24),
  I1 => R1IN_ADD_1(7),
  O => R1IN_ADD_2_AXB_7);
R1IN_ADD_2_AXB_8_Z4576: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(25),
  I1 => R1IN_ADD_1(8),
  O => R1IN_ADD_2_AXB_8);
R1IN_ADD_2_AXB_9_Z4577: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(26),
  I1 => R1IN_ADD_1(9),
  O => R1IN_ADD_2_AXB_9);
R1IN_ADD_2_AXB_10_Z4578: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(27),
  I1 => R1IN_ADD_1(10),
  O => R1IN_ADD_2_AXB_10);
R1IN_ADD_2_AXB_11_Z4579: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(28),
  I1 => R1IN_ADD_1(11),
  O => R1IN_ADD_2_AXB_11);
R1IN_ADD_2_AXB_12_Z4580: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(29),
  I1 => R1IN_ADD_1(12),
  O => R1IN_ADD_2_AXB_12);
R1IN_ADD_2_AXB_13_Z4581: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(30),
  I1 => R1IN_ADD_1(13),
  O => R1IN_ADD_2_AXB_13);
R1IN_ADD_2_AXB_14_Z4582: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(31),
  I1 => R1IN_ADD_1(14),
  O => R1IN_ADD_2_AXB_14);
R1IN_ADD_2_AXB_15_Z4583: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(32),
  I1 => R1IN_ADD_1(15),
  O => R1IN_ADD_2_AXB_15);
R1IN_ADD_2_AXB_16_Z4584: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(33),
  I1 => R1IN_ADD_1(16),
  O => R1IN_ADD_2_AXB_16);
R1IN_ADD_2_AXB_17_Z4585: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(0),
  I1 => R1IN_ADD_1(17),
  O => R1IN_ADD_2_AXB_17);
R1IN_ADD_2_AXB_18_Z4586: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(1),
  I1 => R1IN_ADD_1(18),
  O => R1IN_ADD_2_AXB_18);
R1IN_ADD_2_AXB_19_Z4587: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(2),
  I1 => R1IN_ADD_1(19),
  O => R1IN_ADD_2_AXB_19);
R1IN_ADD_2_AXB_20_Z4588: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(3),
  I1 => R1IN_ADD_1(20),
  O => R1IN_ADD_2_AXB_20);
R1IN_ADD_2_AXB_21_Z4589: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(4),
  I1 => R1IN_ADD_1(21),
  O => R1IN_ADD_2_AXB_21);
R1IN_ADD_2_AXB_22_Z4590: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(5),
  I1 => R1IN_ADD_1(22),
  O => R1IN_ADD_2_AXB_22);
R1IN_ADD_2_AXB_23_Z4591: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(6),
  I1 => R1IN_ADD_1(23),
  O => R1IN_ADD_2_AXB_23);
R1IN_ADD_2_AXB_24_Z4592: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(7),
  I1 => R1IN_ADD_1(24),
  O => R1IN_ADD_2_AXB_24);
R1IN_ADD_2_AXB_25_Z4593: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(8),
  I1 => R1IN_ADD_1(25),
  O => R1IN_ADD_2_AXB_25);
R1IN_ADD_2_AXB_26_Z4594: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(9),
  I1 => R1IN_ADD_1(26),
  O => R1IN_ADD_2_AXB_26);
R1IN_ADD_2_AXB_27_Z4595: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(10),
  I1 => R1IN_ADD_1(27),
  O => R1IN_ADD_2_AXB_27);
R1IN_ADD_2_AXB_28_Z4596: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(11),
  I1 => R1IN_ADD_1(28),
  O => R1IN_ADD_2_AXB_28);
R1IN_ADD_2_AXB_29_Z4597: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(12),
  I1 => R1IN_ADD_1(29),
  O => R1IN_ADD_2_AXB_29);
R1IN_ADD_2_AXB_30_Z4598: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(13),
  I1 => R1IN_ADD_1(30),
  O => R1IN_ADD_2_AXB_30);
R1IN_ADD_2_AXB_31_Z4599: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(14),
  I1 => R1IN_ADD_1(31),
  O => R1IN_ADD_2_AXB_31);
R1IN_ADD_2_AXB_32_Z4600: LUT4 
generic map(
  INIT => X"95A6"
)
port map (
  I0 => R1IN_4FF(15),
  I1 => R1IN_ADD_1_0_CRY_31,
  I2 => R1IN_ADD_1_1_0_AXB_0,
  I3 => R1IN_ADD_1_1_AXB_0,
  O => R1IN_ADD_2_AXB_32);
R1IN_ADD_2_AXB_33_Z4601: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1379,
  I1 => N_1565,
  I2 => R1IN_4FF(16),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_33);
R1IN_ADD_2_AXB_34_Z4602: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1381,
  I1 => N_1566,
  I2 => R1IN_4(17),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_34);
R1IN_ADD_2_AXB_35_Z4603: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1383,
  I1 => N_1567,
  I2 => R1IN_4(18),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_35);
R1IN_ADD_2_AXB_36_Z4604: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1385,
  I1 => N_1568,
  I2 => R1IN_4(19),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_36);
R1IN_ADD_2_AXB_37_Z4605: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1387,
  I1 => N_1569,
  I2 => R1IN_4(20),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_37);
R1IN_ADD_2_AXB_38_Z4606: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1389,
  I1 => N_1570,
  I2 => R1IN_4(21),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_38);
R1IN_ADD_2_AXB_39_Z4607: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1391,
  I1 => N_1571,
  I2 => R1IN_4(22),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_39);
R1IN_ADD_2_AXB_40_Z4608: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1393,
  I1 => N_1572,
  I2 => R1IN_4(23),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_40);
R1IN_ADD_2_AXB_41_Z4609: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1395,
  I1 => N_1573,
  I2 => R1IN_4(24),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_41);
R1IN_ADD_2_AXB_42_Z4610: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1397,
  I1 => N_1574,
  I2 => R1IN_4(25),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_42);
R1IN_ADD_2_AXB_43_Z4611: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1399,
  I1 => N_1575,
  I2 => R1IN_4(26),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_43);
R1IN_ADD_2_AXB_44_Z4612: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1401,
  I1 => N_1576,
  I2 => R1IN_4(27),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_44);
R1IN_ADD_2_AXB_45_Z4613: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1403,
  I1 => N_1577,
  I2 => R1IN_4(28),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_45);
R1IN_ADD_2_AXB_46_Z4614: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1405,
  I1 => N_1578,
  I2 => R1IN_4(29),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_46);
R1IN_ADD_2_AXB_47_Z4615: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1407,
  I1 => N_1579,
  I2 => R1IN_4(30),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_47);
R1IN_ADD_2_AXB_48_Z4616: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1409,
  I1 => N_1580,
  I2 => R1IN_4(31),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_48);
R1IN_ADD_2_AXB_49_Z4617: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1411,
  I1 => N_1581,
  I2 => R1IN_4(32),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_49);
R1IN_ADD_2_AXB_50_Z4618: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1413,
  I1 => N_1582,
  I2 => R1IN_4(33),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_50);
R1IN_ADD_2_AXB_51_Z4619: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1415,
  I1 => N_1583,
  I2 => R1IN_4(34),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_51);
R1IN_ADD_2_AXB_52_Z4620: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1417,
  I1 => N_1584,
  I2 => R1IN_4(35),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_52);
R1IN_ADD_2_AXB_53_Z4621: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1419,
  I1 => N_1585,
  I2 => R1IN_4(36),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_53);
R1IN_ADD_2_AXB_54_Z4622: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1421,
  I1 => N_1586,
  I2 => R1IN_4(37),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_54);
R1IN_ADD_2_AXB_55_Z4623: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1423,
  I1 => N_1587,
  I2 => R1IN_4(38),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_55);
R1IN_ADD_2_AXB_56_Z4624: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1425,
  I1 => N_1588,
  I2 => R1IN_4(39),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_56);
R1IN_ADD_2_AXB_57_Z4625: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1427,
  I1 => N_1589,
  I2 => R1IN_4(40),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_57);
R1IN_ADD_2_AXB_58_Z4626: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1429,
  I1 => N_1590,
  I2 => R1IN_4(41),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_58);
R1IN_ADD_2_AXB_59_Z4627: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1431,
  I1 => N_1591,
  I2 => R1IN_4(42),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_59);
R1IN_ADD_2_AXB_60_Z4628: LUT4 
generic map(
  INIT => X"3C5A"
)
port map (
  I0 => N_1433,
  I1 => N_1592,
  I2 => R1IN_4(43),
  I3 => R1IN_ADD_1_0_CRY_31,
  O => R1IN_ADD_2_AXB_60);
R1IN_ADD_2_AXB_61_Z4629: LUT4 
generic map(
  INIT => X"596A"
)
port map (
  I0 => R1IN_4(44),
  I1 => R1IN_ADD_1_0_CRY_31,
  I2 => R1IN_ADD_1_1_0_CRY_28,
  I3 => R1IN_ADD_1_1_CRY_28,
  O => R1IN_ADD_2_AXB_61);
R1IN_ADD_2_AXB_62_Z4630: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4(45),
  O => R1IN_ADD_2_AXB_62);
R1IN_ADD_2_AXB_63_Z4631: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4(46),
  O => R1IN_ADD_2_AXB_63);
R1IN_ADD_2_AXB_64_Z4632: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4(47),
  O => R1IN_ADD_2_AXB_64);
R1IN_ADD_2_AXB_65_Z4633: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4(48),
  O => R1IN_ADD_2_AXB_65);
R1IN_ADD_2_AXB_66_Z4634: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4(49),
  O => R1IN_ADD_2_AXB_66);
R1IN_ADD_2_AXB_67_Z4635: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4(50),
  O => R1IN_ADD_2_AXB_67);
R1IN_ADD_2_AXB_68_Z4636: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4(51),
  O => R1IN_ADD_2_AXB_68);
R1IN_ADD_2_AXB_69_Z4637: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4(52),
  O => R1IN_ADD_2_AXB_69);
R1IN_ADD_2_AXB_70_Z4638: LUT3 
generic map(
  INIT => X"72"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35,
  I1 => R1IN_4_ADD_2_1_0_AXB_0,
  I2 => R1IN_4_ADD_2_1_AXB_0,
  O => R1IN_ADD_2_AXB_70);
R1IN_ADD_2_AXB_71_Z4639: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1445,
  I1 => N_1523,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_71);
R1IN_ADD_2_AXB_72_Z4640: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1447,
  I1 => N_1524,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_72);
R1IN_ADD_2_AXB_73_Z4641: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1449,
  I1 => N_1525,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_73);
R1IN_ADD_2_AXB_74_Z4642: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1451,
  I1 => N_1526,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_74);
R1IN_ADD_2_AXB_75_Z4643: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1453,
  I1 => N_1527,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_75);
R1IN_ADD_2_AXB_76_Z4644: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1455,
  I1 => N_1528,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_76);
R1IN_ADD_2_AXB_77_Z4645: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1457,
  I1 => N_1529,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_77);
R1IN_ADD_2_AXB_78_Z4646: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1459,
  I1 => N_1530,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_78);
R1IN_ADD_2_AXB_79_Z4647: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1461,
  I1 => N_1531,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_79);
R1IN_ADD_2_AXB_80_Z4648: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1463,
  I1 => N_1532,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_80);
R1IN_ADD_2_AXB_81_Z4649: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1465,
  I1 => N_1533,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_81);
R1IN_ADD_2_AXB_82_Z4650: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1467,
  I1 => N_1534,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_82);
R1IN_ADD_2_AXB_83_Z4651: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1469,
  I1 => N_1535,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_83);
R1IN_ADD_2_AXB_84_Z4652: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1471,
  I1 => N_1536,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_84);
R1IN_ADD_2_AXB_85_Z4653: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1473,
  I1 => N_1537,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_85);
R1IN_ADD_2_AXB_86_Z4654: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1475,
  I1 => N_1538,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_86);
R1IN_ADD_2_AXB_87_Z4655: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1477,
  I1 => N_1539,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_87);
R1IN_ADD_2_AXB_88_Z4656: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1479,
  I1 => N_1540,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_88);
R1IN_ADD_2_AXB_89_Z4657: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1481,
  I1 => N_1541,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_89);
R1IN_ADD_2_AXB_90_Z4658: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1483,
  I1 => N_1542,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_90);
R1IN_ADD_2_AXB_91_Z4659: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1485,
  I1 => N_1543,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_91);
R1IN_ADD_2_AXB_92_Z4660: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1487,
  I1 => N_1544,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_92);
R1IN_ADD_2_AXB_93_Z4661: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1489,
  I1 => N_1545,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_93);
R1IN_ADD_2_AXB_94_Z4662: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1491,
  I1 => N_1546,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_94);
R1IN_ADD_2_AXB_95_Z4663: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1493,
  I1 => N_1547,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_95);
R1IN_ADD_2_AXB_96_Z4664: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1495,
  I1 => N_1548,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_96);
R1IN_ADD_2_AXB_97_Z4665: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1497,
  I1 => N_1549,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_97);
R1IN_ADD_2_AXB_98_Z4666: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1499,
  I1 => N_1550,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_98);
R1IN_ADD_2_AXB_99_Z4667: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1501,
  I1 => N_1551,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_99);
R1IN_ADD_2_AXB_100_Z4668: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1503,
  I1 => N_1552,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_100);
R1IN_ADD_2_AXB_101_Z4669: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1505,
  I1 => N_1553,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_101);
R1IN_ADD_2_AXB_102_Z4670: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1507,
  I1 => N_1554,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_102);
R1IN_ADD_2_AXB_103_Z4671: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1509,
  I1 => N_1555,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_103);
R1IN_2_ADD_1_AXB_1_Z4672: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F_RETO(18),
  I1 => R1IN_2_2F_RETO(1),
  O => R1IN_2_ADD_1_AXB_1);
R1IN_2_ADD_1_AXB_2_Z4673: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F_RETO(19),
  I1 => R1IN_2_2F_RETO(2),
  O => R1IN_2_ADD_1_AXB_2);
R1IN_2_ADD_1_AXB_3_Z4674: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F_RETO(20),
  I1 => R1IN_2_2F_RETO(3),
  O => R1IN_2_ADD_1_AXB_3);
R1IN_2_ADD_1_AXB_4_Z4675: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F_RETO(21),
  I1 => R1IN_2_2F_RETO(4),
  O => R1IN_2_ADD_1_AXB_4);
R1IN_2_ADD_1_AXB_5_Z4676: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F_RETO(22),
  I1 => R1IN_2_2F_RETO(5),
  O => R1IN_2_ADD_1_AXB_5);
R1IN_2_ADD_1_AXB_6_Z4677: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F_RETO(23),
  I1 => R1IN_2_2F_RETO(6),
  O => R1IN_2_ADD_1_AXB_6);
R1IN_2_ADD_1_AXB_7_Z4678: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F_RETO(24),
  I1 => R1IN_2_2F_RETO(7),
  O => R1IN_2_ADD_1_AXB_7);
R1IN_2_ADD_1_AXB_8_Z4679: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F_RETO(25),
  I1 => R1IN_2_2F_RETO(8),
  O => R1IN_2_ADD_1_AXB_8);
R1IN_2_ADD_1_AXB_9_Z4680: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F_RETO(26),
  I1 => R1IN_2_2F_RETO(9),
  O => R1IN_2_ADD_1_AXB_9);
R1IN_2_ADD_1_AXB_10_Z4681: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F_RETO(27),
  I1 => R1IN_2_2F_RETO(10),
  O => R1IN_2_ADD_1_AXB_10);
R1IN_2_ADD_1_AXB_11_Z4682: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F_RETO(28),
  I1 => R1IN_2_2F_RETO(11),
  O => R1IN_2_ADD_1_AXB_11);
R1IN_2_ADD_1_AXB_12_Z4683: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F_RETO(29),
  I1 => R1IN_2_2F_RETO(12),
  O => R1IN_2_ADD_1_AXB_12);
R1IN_2_ADD_1_AXB_13_Z4684: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F_RETO(30),
  I1 => R1IN_2_2F_RETO(13),
  O => R1IN_2_ADD_1_AXB_13);
R1IN_2_ADD_1_AXB_14_Z4685: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F_RETO(31),
  I1 => R1IN_2_2F_RETO(14),
  O => R1IN_2_ADD_1_AXB_14);
R1IN_2_ADD_1_AXB_15_Z4686: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F_RETO(32),
  I1 => R1IN_2_2F_RETO(15),
  O => R1IN_2_ADD_1_AXB_15);
R1IN_2_ADD_1_AXB_16_Z4687: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F_RETO(33),
  I1 => R1IN_2_2F_RETO(16),
  O => R1IN_2_ADD_1_AXB_16);
R1IN_2_ADD_1_AXB_17_Z4688: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(17),
  O => R1IN_2_ADD_1_AXB_17);
R1IN_2_ADD_1_AXB_18_Z4689: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(18),
  O => R1IN_2_ADD_1_AXB_18);
R1IN_2_ADD_1_AXB_19_Z4690: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(19),
  O => R1IN_2_ADD_1_AXB_19);
R1IN_2_ADD_1_AXB_20_Z4691: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(20),
  O => R1IN_2_ADD_1_AXB_20);
R1IN_2_ADD_1_AXB_21_Z4692: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(21),
  O => R1IN_2_ADD_1_AXB_21);
R1IN_2_ADD_1_AXB_22_Z4693: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(22),
  O => R1IN_2_ADD_1_AXB_22);
R1IN_2_ADD_1_AXB_23_Z4694: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(23),
  O => R1IN_2_ADD_1_AXB_23);
R1IN_2_ADD_1_AXB_24_Z4695: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(24),
  O => R1IN_2_ADD_1_AXB_24);
R1IN_2_ADD_1_AXB_25_Z4696: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(25),
  O => R1IN_2_ADD_1_AXB_25);
R1IN_2_ADD_1_AXB_26_Z4697: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(26),
  O => R1IN_2_ADD_1_AXB_26);
R1IN_2_ADD_1_AXB_27_Z4698: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(27),
  O => R1IN_2_ADD_1_AXB_27);
R1IN_2_ADD_1_AXB_28_Z4699: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(28),
  O => R1IN_2_ADD_1_AXB_28);
R1IN_2_ADD_1_AXB_29_Z4700: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(29),
  O => R1IN_2_ADD_1_AXB_29);
R1IN_2_ADD_1_AXB_30_Z4701: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(30),
  O => R1IN_2_ADD_1_AXB_30);
R1IN_2_ADD_1_AXB_31_Z4702: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(31),
  O => R1IN_2_ADD_1_AXB_31);
R1IN_2_ADD_1_AXB_32_Z4703: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(32),
  O => R1IN_2_ADD_1_AXB_32);
R1IN_2_ADD_1_AXB_33_Z4704: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(33),
  O => R1IN_2_ADD_1_AXB_33);
R1IN_2_ADD_1_AXB_34_Z4705: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(34),
  O => R1IN_2_ADD_1_AXB_34);
R1IN_2_ADD_1_AXB_35_Z4706: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(35),
  O => R1IN_2_ADD_1_AXB_35);
R1IN_2_ADD_1_AXB_36_Z4707: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(36),
  O => R1IN_2_ADD_1_AXB_36);
R1IN_2_ADD_1_AXB_37_Z4708: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(37),
  O => R1IN_2_ADD_1_AXB_37);
R1IN_2_ADD_1_AXB_38_Z4709: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(38),
  O => R1IN_2_ADD_1_AXB_38);
R1IN_2_ADD_1_AXB_39_Z4710: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(39),
  O => R1IN_2_ADD_1_AXB_39);
R1IN_2_ADD_1_AXB_40_Z4711: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(40),
  O => R1IN_2_ADD_1_AXB_40);
R1IN_2_ADD_1_AXB_41_Z4712: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(41),
  O => R1IN_2_ADD_1_AXB_41);
R1IN_2_ADD_1_AXB_42_Z4713: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(42),
  O => R1IN_2_ADD_1_AXB_42);
R1IN_4_ADD_1_AXB_1_Z4714: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(1),
  I1 => R1IN_4_3F_RETO(1),
  O => R1IN_4_ADD_1_AXB_1);
R1IN_4_ADD_1_AXB_2_Z4715: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(2),
  I1 => R1IN_4_3F_RETO(2),
  O => R1IN_4_ADD_1_AXB_2);
R1IN_4_ADD_1_AXB_3_Z4716: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(3),
  I1 => R1IN_4_3F_RETO(3),
  O => R1IN_4_ADD_1_AXB_3);
R1IN_4_ADD_1_AXB_4_Z4717: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(4),
  I1 => R1IN_4_3F_RETO(4),
  O => R1IN_4_ADD_1_AXB_4);
R1IN_4_ADD_1_AXB_5_Z4718: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(5),
  I1 => R1IN_4_3F_RETO(5),
  O => R1IN_4_ADD_1_AXB_5);
R1IN_4_ADD_1_AXB_6_Z4719: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(6),
  I1 => R1IN_4_3F_RETO(6),
  O => R1IN_4_ADD_1_AXB_6);
R1IN_4_ADD_1_AXB_7_Z4720: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(7),
  I1 => R1IN_4_3F_RETO(7),
  O => R1IN_4_ADD_1_AXB_7);
R1IN_4_ADD_1_AXB_8_Z4721: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(8),
  I1 => R1IN_4_3F_RETO(8),
  O => R1IN_4_ADD_1_AXB_8);
R1IN_4_ADD_1_AXB_9_Z4722: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(9),
  I1 => R1IN_4_3F_RETO(9),
  O => R1IN_4_ADD_1_AXB_9);
R1IN_4_ADD_1_AXB_10_Z4723: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(10),
  I1 => R1IN_4_3F_RETO(10),
  O => R1IN_4_ADD_1_AXB_10);
R1IN_4_ADD_1_AXB_11_Z4724: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(11),
  I1 => R1IN_4_3F_RETO(11),
  O => R1IN_4_ADD_1_AXB_11);
R1IN_4_ADD_1_AXB_12_Z4725: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(12),
  I1 => R1IN_4_3F_RETO(12),
  O => R1IN_4_ADD_1_AXB_12);
R1IN_4_ADD_1_AXB_13_Z4726: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(13),
  I1 => R1IN_4_3F_RETO(13),
  O => R1IN_4_ADD_1_AXB_13);
R1IN_4_ADD_1_AXB_14_Z4727: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(14),
  I1 => R1IN_4_3F_RETO(14),
  O => R1IN_4_ADD_1_AXB_14);
R1IN_4_ADD_1_AXB_15_Z4728: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(15),
  I1 => R1IN_4_3F_RETO(15),
  O => R1IN_4_ADD_1_AXB_15);
R1IN_4_ADD_1_AXB_16_Z4729: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(16),
  I1 => R1IN_4_3F_RETO(16),
  O => R1IN_4_ADD_1_AXB_16);
R1IN_4_ADD_1_AXB_17_Z4730: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(17),
  I1 => R1IN_4_3F_RETO(17),
  O => R1IN_4_ADD_1_AXB_17);
R1IN_4_ADD_1_AXB_18_Z4731: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(18),
  I1 => R1IN_4_3F_RETO(18),
  O => R1IN_4_ADD_1_AXB_18);
R1IN_4_ADD_1_AXB_19_Z4732: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(19),
  I1 => R1IN_4_3F_RETO(19),
  O => R1IN_4_ADD_1_AXB_19);
R1IN_4_ADD_1_AXB_20_Z4733: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(20),
  I1 => R1IN_4_3F_RETO(20),
  O => R1IN_4_ADD_1_AXB_20);
R1IN_4_ADD_1_AXB_21_Z4734: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(21),
  I1 => R1IN_4_3F_RETO(21),
  O => R1IN_4_ADD_1_AXB_21);
R1IN_4_ADD_1_AXB_22_Z4735: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(22),
  I1 => R1IN_4_3F_RETO(22),
  O => R1IN_4_ADD_1_AXB_22);
R1IN_4_ADD_1_AXB_23_Z4736: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(23),
  I1 => R1IN_4_3F_RETO(23),
  O => R1IN_4_ADD_1_AXB_23);
R1IN_4_ADD_1_AXB_24_Z4737: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(24),
  I1 => R1IN_4_3F_RETO(24),
  O => R1IN_4_ADD_1_AXB_24);
R1IN_4_ADD_1_AXB_25_Z4738: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(25),
  I1 => R1IN_4_3F_RETO(25),
  O => R1IN_4_ADD_1_AXB_25);
R1IN_4_ADD_1_AXB_26_Z4739: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(26),
  I1 => R1IN_4_3F_RETO(26),
  O => R1IN_4_ADD_1_AXB_26);
R1IN_4_ADD_1_AXB_27_Z4740: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(27),
  I1 => R1IN_4_3F_RETO(27),
  O => R1IN_4_ADD_1_AXB_27);
R1IN_4_ADD_1_AXB_28_Z4741: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(28),
  I1 => R1IN_4_3F_RETO(28),
  O => R1IN_4_ADD_1_AXB_28);
R1IN_4_ADD_1_AXB_29_Z4742: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(29),
  I1 => R1IN_4_3F_RETO(29),
  O => R1IN_4_ADD_1_AXB_29);
R1IN_4_ADD_1_AXB_30_Z4743: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(30),
  I1 => R1IN_4_3F_RETO(30),
  O => R1IN_4_ADD_1_AXB_30);
R1IN_4_ADD_1_AXB_31_Z4744: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(31),
  I1 => R1IN_4_3F_RETO(31),
  O => R1IN_4_ADD_1_AXB_31);
R1IN_4_ADD_1_AXB_32_Z4745: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(32),
  I1 => R1IN_4_3F_RETO(32),
  O => R1IN_4_ADD_1_AXB_32);
R1IN_4_ADD_1_AXB_33_Z4746: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(33),
  I1 => R1IN_4_3F_RETO(33),
  O => R1IN_4_ADD_1_AXB_33);
R1IN_4_ADD_1_AXB_34_Z4747: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(34),
  I1 => R1IN_4_3F_RETO(34),
  O => R1IN_4_ADD_1_AXB_34);
R1IN_4_ADD_1_AXB_35_Z4748: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(35),
  I1 => R1IN_4_3F_RETO(35),
  O => R1IN_4_ADD_1_AXB_35);
R1IN_4_ADD_1_AXB_36_Z4749: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(36),
  I1 => R1IN_4_3F_RETO(36),
  O => R1IN_4_ADD_1_AXB_36);
R1IN_4_ADD_1_AXB_37_Z4750: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(37),
  I1 => R1IN_4_3F_RETO(37),
  O => R1IN_4_ADD_1_AXB_37);
R1IN_4_ADD_1_AXB_38_Z4751: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(38),
  I1 => R1IN_4_3F_RETO(38),
  O => R1IN_4_ADD_1_AXB_38);
R1IN_4_ADD_1_AXB_39_Z4752: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(39),
  I1 => R1IN_4_3F_RETO(39),
  O => R1IN_4_ADD_1_AXB_39);
R1IN_4_ADD_1_AXB_40_Z4753: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(40),
  I1 => R1IN_4_3F_RETO(40),
  O => R1IN_4_ADD_1_AXB_40);
R1IN_4_ADD_1_AXB_41_Z4754: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(41),
  I1 => R1IN_4_3F_RETO(41),
  O => R1IN_4_ADD_1_AXB_41);
R1IN_4_ADD_1_AXB_42_Z4755: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(42),
  I1 => R1IN_4_3F_RETO(42),
  O => R1IN_4_ADD_1_AXB_42);
R1IN_4_ADD_1_AXB_43_Z4756: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F_RETO(43),
  I1 => R1IN_4_3F_RETO(43),
  O => R1IN_4_ADD_1_AXB_43);
R1IN_ADD_1_1_AXB_28_Z4757: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(60),
  I1 => R1IN_3(60),
  O => R1IN_ADD_1_1_AXB_28);
R1_PIPE_34: FDE port map (
    Q => R1IN_4_ADD_1,
    D => R1IN_4_2(0),
    C => CLK,
    CE => EN);
R1_PIPE_283: FDE port map (
    Q => R1IN_4_2F(1),
    D => R1IN_4_2(1),
    C => CLK,
    CE => EN);
R1_PIPE_284: FDE port map (
    Q => R1IN_4_2F(2),
    D => R1IN_4_2(2),
    C => CLK,
    CE => EN);
R1_PIPE_285: FDE port map (
    Q => R1IN_4_2F(3),
    D => R1IN_4_2(3),
    C => CLK,
    CE => EN);
R1_PIPE_286: FDE port map (
    Q => R1IN_4_2F(4),
    D => R1IN_4_2(4),
    C => CLK,
    CE => EN);
R1_PIPE_287: FDE port map (
    Q => R1IN_4_2F(5),
    D => R1IN_4_2(5),
    C => CLK,
    CE => EN);
R1_PIPE_288: FDE port map (
    Q => R1IN_4_2F(6),
    D => R1IN_4_2(6),
    C => CLK,
    CE => EN);
R1_PIPE_289: FDE port map (
    Q => R1IN_4_2F(7),
    D => R1IN_4_2(7),
    C => CLK,
    CE => EN);
R1_PIPE_290: FDE port map (
    Q => R1IN_4_2F(8),
    D => R1IN_4_2(8),
    C => CLK,
    CE => EN);
R1_PIPE_291: FDE port map (
    Q => R1IN_4_2F(9),
    D => R1IN_4_2(9),
    C => CLK,
    CE => EN);
R1_PIPE_292: FDE port map (
    Q => R1IN_4_2F(10),
    D => R1IN_4_2(10),
    C => CLK,
    CE => EN);
R1_PIPE_293: FDE port map (
    Q => R1IN_4_2F(11),
    D => R1IN_4_2(11),
    C => CLK,
    CE => EN);
R1_PIPE_294: FDE port map (
    Q => R1IN_4_2F(12),
    D => R1IN_4_2(12),
    C => CLK,
    CE => EN);
R1_PIPE_295: FDE port map (
    Q => R1IN_4_2F(13),
    D => R1IN_4_2(13),
    C => CLK,
    CE => EN);
R1_PIPE_296: FDE port map (
    Q => R1IN_4_2F(14),
    D => R1IN_4_2(14),
    C => CLK,
    CE => EN);
R1_PIPE_297: FDE port map (
    Q => R1IN_4_2F(15),
    D => R1IN_4_2(15),
    C => CLK,
    CE => EN);
R1_PIPE_298: FDE port map (
    Q => R1IN_4_2F(16),
    D => R1IN_4_2(16),
    C => CLK,
    CE => EN);
R1_PIPE_326: FDE port map (
    Q => R1IN_4_3F(0),
    D => R1IN_4_3(0),
    C => CLK,
    CE => EN);
R1_PIPE_327: FDE port map (
    Q => R1IN_4_3F(1),
    D => R1IN_4_3(1),
    C => CLK,
    CE => EN);
R1_PIPE_328: FDE port map (
    Q => R1IN_4_3F(2),
    D => R1IN_4_3(2),
    C => CLK,
    CE => EN);
R1_PIPE_329: FDE port map (
    Q => R1IN_4_3F(3),
    D => R1IN_4_3(3),
    C => CLK,
    CE => EN);
R1_PIPE_330: FDE port map (
    Q => R1IN_4_3F(4),
    D => R1IN_4_3(4),
    C => CLK,
    CE => EN);
R1_PIPE_331: FDE port map (
    Q => R1IN_4_3F(5),
    D => R1IN_4_3(5),
    C => CLK,
    CE => EN);
R1_PIPE_332: FDE port map (
    Q => R1IN_4_3F(6),
    D => R1IN_4_3(6),
    C => CLK,
    CE => EN);
R1_PIPE_333: FDE port map (
    Q => R1IN_4_3F(7),
    D => R1IN_4_3(7),
    C => CLK,
    CE => EN);
R1_PIPE_334: FDE port map (
    Q => R1IN_4_3F(8),
    D => R1IN_4_3(8),
    C => CLK,
    CE => EN);
R1_PIPE_335: FDE port map (
    Q => R1IN_4_3F(9),
    D => R1IN_4_3(9),
    C => CLK,
    CE => EN);
R1_PIPE_336: FDE port map (
    Q => R1IN_4_3F(10),
    D => R1IN_4_3(10),
    C => CLK,
    CE => EN);
R1_PIPE_337: FDE port map (
    Q => R1IN_4_3F(11),
    D => R1IN_4_3(11),
    C => CLK,
    CE => EN);
R1_PIPE_338: FDE port map (
    Q => R1IN_4_3F(12),
    D => R1IN_4_3(12),
    C => CLK,
    CE => EN);
R1_PIPE_339: FDE port map (
    Q => R1IN_4_3F(13),
    D => R1IN_4_3(13),
    C => CLK,
    CE => EN);
R1_PIPE_340: FDE port map (
    Q => R1IN_4_3F(14),
    D => R1IN_4_3(14),
    C => CLK,
    CE => EN);
R1_PIPE_341: FDE port map (
    Q => R1IN_4_3F(15),
    D => R1IN_4_3(15),
    C => CLK,
    CE => EN);
R1_PIPE_342: FDE port map (
    Q => R1IN_4_3F(16),
    D => R1IN_4_3(16),
    C => CLK,
    CE => EN);
R1_PIPE_105: FDE port map (
    Q => R1IN_2_ADD_1,
    D => R1IN_2_2(0),
    C => CLK,
    CE => EN);
R1_PIPE_589: FDE port map (
    Q => R1IN_2_2F(1),
    D => R1IN_2_2(1),
    C => CLK,
    CE => EN);
R1_PIPE_590: FDE port map (
    Q => R1IN_2_2F(2),
    D => R1IN_2_2(2),
    C => CLK,
    CE => EN);
R1_PIPE_591: FDE port map (
    Q => R1IN_2_2F(3),
    D => R1IN_2_2(3),
    C => CLK,
    CE => EN);
R1_PIPE_592: FDE port map (
    Q => R1IN_2_2F(4),
    D => R1IN_2_2(4),
    C => CLK,
    CE => EN);
R1_PIPE_593: FDE port map (
    Q => R1IN_2_2F(5),
    D => R1IN_2_2(5),
    C => CLK,
    CE => EN);
R1_PIPE_594: FDE port map (
    Q => R1IN_2_2F(6),
    D => R1IN_2_2(6),
    C => CLK,
    CE => EN);
R1_PIPE_595: FDE port map (
    Q => R1IN_2_2F(7),
    D => R1IN_2_2(7),
    C => CLK,
    CE => EN);
R1_PIPE_596: FDE port map (
    Q => R1IN_2_2F(8),
    D => R1IN_2_2(8),
    C => CLK,
    CE => EN);
R1_PIPE_597: FDE port map (
    Q => R1IN_2_2F(9),
    D => R1IN_2_2(9),
    C => CLK,
    CE => EN);
R1_PIPE_598: FDE port map (
    Q => R1IN_2_2F(10),
    D => R1IN_2_2(10),
    C => CLK,
    CE => EN);
R1_PIPE_599: FDE port map (
    Q => R1IN_2_2F(11),
    D => R1IN_2_2(11),
    C => CLK,
    CE => EN);
R1_PIPE_600: FDE port map (
    Q => R1IN_2_2F(12),
    D => R1IN_2_2(12),
    C => CLK,
    CE => EN);
R1_PIPE_601: FDE port map (
    Q => R1IN_2_2F(13),
    D => R1IN_2_2(13),
    C => CLK,
    CE => EN);
R1_PIPE_602: FDE port map (
    Q => R1IN_2_2F(14),
    D => R1IN_2_2(14),
    C => CLK,
    CE => EN);
R1_PIPE_603: FDE port map (
    Q => R1IN_2_2F(15),
    D => R1IN_2_2(15),
    C => CLK,
    CE => EN);
R1_PIPE_604: FDE port map (
    Q => R1IN_2_2F(16),
    D => R1IN_2_2(16),
    C => CLK,
    CE => EN);
R1_PIPE_484: FDE port map (
    Q => R1IN_3_ADD_1,
    D => R1IN_3_2(0),
    C => CLK,
    CE => EN);
R1_PIPE_649: FDE port map (
    Q => R1IN_3_2F(1),
    D => R1IN_3_2(1),
    C => CLK,
    CE => EN);
R1_PIPE_650: FDE port map (
    Q => R1IN_3_2F(2),
    D => R1IN_3_2(2),
    C => CLK,
    CE => EN);
R1_PIPE_651: FDE port map (
    Q => R1IN_3_2F(3),
    D => R1IN_3_2(3),
    C => CLK,
    CE => EN);
R1_PIPE_652: FDE port map (
    Q => R1IN_3_2F(4),
    D => R1IN_3_2(4),
    C => CLK,
    CE => EN);
R1_PIPE_653: FDE port map (
    Q => R1IN_3_2F(5),
    D => R1IN_3_2(5),
    C => CLK,
    CE => EN);
R1_PIPE_654: FDE port map (
    Q => R1IN_3_2F(6),
    D => R1IN_3_2(6),
    C => CLK,
    CE => EN);
R1_PIPE_655: FDE port map (
    Q => R1IN_3_2F(7),
    D => R1IN_3_2(7),
    C => CLK,
    CE => EN);
R1_PIPE_656: FDE port map (
    Q => R1IN_3_2F(8),
    D => R1IN_3_2(8),
    C => CLK,
    CE => EN);
R1_PIPE_657: FDE port map (
    Q => R1IN_3_2F(9),
    D => R1IN_3_2(9),
    C => CLK,
    CE => EN);
R1_PIPE_658: FDE port map (
    Q => R1IN_3_2F(10),
    D => R1IN_3_2(10),
    C => CLK,
    CE => EN);
R1_PIPE_659: FDE port map (
    Q => R1IN_3_2F(11),
    D => R1IN_3_2(11),
    C => CLK,
    CE => EN);
R1_PIPE_660: FDE port map (
    Q => R1IN_3_2F(12),
    D => R1IN_3_2(12),
    C => CLK,
    CE => EN);
R1_PIPE_661: FDE port map (
    Q => R1IN_3_2F(13),
    D => R1IN_3_2(13),
    C => CLK,
    CE => EN);
R1_PIPE_662: FDE port map (
    Q => R1IN_3_2F(14),
    D => R1IN_3_2(14),
    C => CLK,
    CE => EN);
R1_PIPE_663: FDE port map (
    Q => R1IN_3_2F(15),
    D => R1IN_3_2(15),
    C => CLK,
    CE => EN);
R1_PIPE_664: FDE port map (
    Q => R1IN_3_2F(16),
    D => R1IN_3_2(16),
    C => CLK,
    CE => EN);
R2_PIPE_136_RET_1: FDE port map (
    Q => R1IN_3F_RETO(0),
    D => R1IN_3F(0),
    C => CLK,
    CE => EN);
R2_PIPE_136_RET_3: FDE port map (
    Q => R1IN_3F_RETO(1),
    D => R1IN_3F(1),
    C => CLK,
    CE => EN);
R2_PIPE_136_RET_5: FDE port map (
    Q => R1IN_3F_RETO(2),
    D => R1IN_3F(2),
    C => CLK,
    CE => EN);
R2_PIPE_136_RET_7: FDE port map (
    Q => R1IN_3F_RETO(3),
    D => R1IN_3F(3),
    C => CLK,
    CE => EN);
R2_PIPE_136_RET_9: FDE port map (
    Q => R1IN_3F_RETO(4),
    D => R1IN_3F(4),
    C => CLK,
    CE => EN);
R2_PIPE_136_RET_11: FDE port map (
    Q => R1IN_3F_RETO(5),
    D => R1IN_3F(5),
    C => CLK,
    CE => EN);
R2_PIPE_136_RET_13: FDE port map (
    Q => R1IN_3F_RETO(6),
    D => R1IN_3F(6),
    C => CLK,
    CE => EN);
R2_PIPE_136_RET_15: FDE port map (
    Q => R1IN_3F_RETO(7),
    D => R1IN_3F(7),
    C => CLK,
    CE => EN);
R2_PIPE_136_RET_17: FDE port map (
    Q => R1IN_3F_RETO(8),
    D => R1IN_3F(8),
    C => CLK,
    CE => EN);
R2_PIPE_136_RET_19: FDE port map (
    Q => R1IN_3F_RETO(9),
    D => R1IN_3F(9),
    C => CLK,
    CE => EN);
R2_PIPE_136_RET_21: FDE port map (
    Q => R1IN_3F_RETO(10),
    D => R1IN_3F(10),
    C => CLK,
    CE => EN);
R2_PIPE_136_RET_23: FDE port map (
    Q => R1IN_3F_RETO(11),
    D => R1IN_3F(11),
    C => CLK,
    CE => EN);
R2_PIPE_136_RET_25: FDE port map (
    Q => R1IN_3F_RETO(12),
    D => R1IN_3F(12),
    C => CLK,
    CE => EN);
R2_PIPE_136_RET_27: FDE port map (
    Q => R1IN_3F_RETO(13),
    D => R1IN_3F(13),
    C => CLK,
    CE => EN);
R2_PIPE_136_RET_29: FDE port map (
    Q => R1IN_3F_RETO(14),
    D => R1IN_3F(14),
    C => CLK,
    CE => EN);
R2_PIPE_136_RET_31: FDE port map (
    Q => R1IN_3F_RETO(15),
    D => R1IN_3F(15),
    C => CLK,
    CE => EN);
R2_PIPE_136_RET_33: FDE port map (
    Q => R1IN_3F_RETO(16),
    D => R1IN_3F(16),
    C => CLK,
    CE => EN);
R2_PIPE_136_RET_35: FDE port map (
    Q => R1IN_3_1F_RETO(17),
    D => R1IN_3_1F(17),
    C => CLK,
    CE => EN);
R2_PIPE_136_RET_36: FDE port map (
    Q => R1IN_3_ADD_1_RETO,
    D => R1IN_3_ADD_1,
    C => CLK,
    CE => EN);
R2_PIPE_69_RET_34: FDE port map (
    Q => R1IN_4_4F_RETO(0),
    D => R1IN_4_4F(0),
    C => CLK,
    CE => EN);
R2_PIPE_69_RET_36: FDE port map (
    Q => R1IN_4_4F_RETO(1),
    D => R1IN_4_4F(1),
    C => CLK,
    CE => EN);
R2_PIPE_69_RET_38: FDE port map (
    Q => R1IN_4_4F_RETO(2),
    D => R1IN_4_4F(2),
    C => CLK,
    CE => EN);
R2_PIPE_69_RET_40: FDE port map (
    Q => R1IN_4_4F_RETO(3),
    D => R1IN_4_4F(3),
    C => CLK,
    CE => EN);
R2_PIPE_69_RET_42: FDE port map (
    Q => R1IN_4_4F_RETO(4),
    D => R1IN_4_4F(4),
    C => CLK,
    CE => EN);
R2_PIPE_69_RET_44: FDE port map (
    Q => R1IN_4_4F_RETO(5),
    D => R1IN_4_4F(5),
    C => CLK,
    CE => EN);
R2_PIPE_69_RET_46: FDE port map (
    Q => R1IN_4_4F_RETO(6),
    D => R1IN_4_4F(6),
    C => CLK,
    CE => EN);
R2_PIPE_69_RET_48: FDE port map (
    Q => R1IN_4_4F_RETO(7),
    D => R1IN_4_4F(7),
    C => CLK,
    CE => EN);
R2_PIPE_69_RET_50: FDE port map (
    Q => R1IN_4_4F_RETO(8),
    D => R1IN_4_4F(8),
    C => CLK,
    CE => EN);
R2_PIPE_69_RET_52: FDE port map (
    Q => R1IN_4_4F_RETO(9),
    D => R1IN_4_4F(9),
    C => CLK,
    CE => EN);
R2_PIPE_69_RET_54: FDE port map (
    Q => R1IN_4_4F_RETO(10),
    D => R1IN_4_4F(10),
    C => CLK,
    CE => EN);
R2_PIPE_69_RET_56: FDE port map (
    Q => R1IN_4_4F_RETO(11),
    D => R1IN_4_4F(11),
    C => CLK,
    CE => EN);
R2_PIPE_69_RET_58: FDE port map (
    Q => R1IN_4_4F_RETO(12),
    D => R1IN_4_4F(12),
    C => CLK,
    CE => EN);
R2_PIPE_69_RET_60: FDE port map (
    Q => R1IN_4_4F_RETO(13),
    D => R1IN_4_4F(13),
    C => CLK,
    CE => EN);
R2_PIPE_69_RET_62: FDE port map (
    Q => R1IN_4_4F_RETO(14),
    D => R1IN_4_4F(14),
    C => CLK,
    CE => EN);
R2_PIPE_69_RET_64: FDE port map (
    Q => R1IN_4_4F_RETO(15),
    D => R1IN_4_4F(15),
    C => CLK,
    CE => EN);
R2_PIPE_69_RET_66: FDE port map (
    Q => R1IN_4_4F_RETO(16),
    D => R1IN_4_4F(16),
    C => CLK,
    CE => EN);
R2_PIPE_69_RET_68: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(0),
    D => R1IN_4_4_ADD_1F(0),
    C => CLK,
    CE => EN);
R2_PIPE_69_RET_69: FDE port map (
    Q => R1IN_4_4_ADD_2_RETO,
    D => R1IN_4_4_ADD_2,
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_119: FDE port map (
    Q => R1IN_3_1F_RETO_0(17),
    D => R1IN_3_1F(17),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_120: FDE port map (
    Q => R1IN_3_ADD_1_RETO_0,
    D => R1IN_3_ADD_1,
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_121: FDE port map (
    Q => R1IN_3_1F_RETO(18),
    D => R1IN_3_1F(18),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_122: FDE port map (
    Q => R1IN_3_2F_RETO(1),
    D => R1IN_3_2F(1),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_123: FDE port map (
    Q => R1IN_3_1F_RETO(19),
    D => R1IN_3_1F(19),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_124: FDE port map (
    Q => R1IN_3_2F_RETO(2),
    D => R1IN_3_2F(2),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_125: FDE port map (
    Q => R1IN_3_1F_RETO(20),
    D => R1IN_3_1F(20),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_126: FDE port map (
    Q => R1IN_3_2F_RETO(3),
    D => R1IN_3_2F(3),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_127: FDE port map (
    Q => R1IN_3_1F_RETO(21),
    D => R1IN_3_1F(21),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_128: FDE port map (
    Q => R1IN_3_2F_RETO(4),
    D => R1IN_3_2F(4),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_129: FDE port map (
    Q => R1IN_3_1F_RETO(22),
    D => R1IN_3_1F(22),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_130: FDE port map (
    Q => R1IN_3_2F_RETO(5),
    D => R1IN_3_2F(5),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_131: FDE port map (
    Q => R1IN_3_1F_RETO(23),
    D => R1IN_3_1F(23),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_132: FDE port map (
    Q => R1IN_3_2F_RETO(6),
    D => R1IN_3_2F(6),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_133: FDE port map (
    Q => R1IN_3_1F_RETO(24),
    D => R1IN_3_1F(24),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_134: FDE port map (
    Q => R1IN_3_2F_RETO(7),
    D => R1IN_3_2F(7),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_135: FDE port map (
    Q => R1IN_3_1F_RETO(25),
    D => R1IN_3_1F(25),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_136: FDE port map (
    Q => R1IN_3_2F_RETO(8),
    D => R1IN_3_2F(8),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_137: FDE port map (
    Q => R1IN_3_1F_RETO(26),
    D => R1IN_3_1F(26),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_138: FDE port map (
    Q => R1IN_3_2F_RETO(9),
    D => R1IN_3_2F(9),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_139: FDE port map (
    Q => R1IN_3_1F_RETO(27),
    D => R1IN_3_1F(27),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_140: FDE port map (
    Q => R1IN_3_2F_RETO(10),
    D => R1IN_3_2F(10),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_141: FDE port map (
    Q => R1IN_3_1F_RETO(28),
    D => R1IN_3_1F(28),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_142: FDE port map (
    Q => R1IN_3_2F_RETO(11),
    D => R1IN_3_2F(11),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_143: FDE port map (
    Q => R1IN_3_1F_RETO(29),
    D => R1IN_3_1F(29),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_144: FDE port map (
    Q => R1IN_3_2F_RETO(12),
    D => R1IN_3_2F(12),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_145: FDE port map (
    Q => R1IN_3_1F_RETO(30),
    D => R1IN_3_1F(30),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_146: FDE port map (
    Q => R1IN_3_2F_RETO(13),
    D => R1IN_3_2F(13),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_147: FDE port map (
    Q => R1IN_3_1F_RETO(31),
    D => R1IN_3_1F(31),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_148: FDE port map (
    Q => R1IN_3_2F_RETO(14),
    D => R1IN_3_2F(14),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_149: FDE port map (
    Q => R1IN_3_1F_RETO(32),
    D => R1IN_3_1F(32),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_150: FDE port map (
    Q => R1IN_3_2F_RETO(15),
    D => R1IN_3_2F(15),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_151: FDE port map (
    Q => R1IN_3_1F_RETO(33),
    D => R1IN_3_1F(33),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_152: FDE port map (
    Q => R1IN_3_2F_RETO(16),
    D => R1IN_3_2F(16),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_153: FDE port map (
    Q => R1IN_3_2F_RETO(17),
    D => R1IN_3_2F(17),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_154: FDE port map (
    Q => R1IN_3_2F_RETO(18),
    D => R1IN_3_2F(18),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_155: FDE port map (
    Q => R1IN_3_2F_RETO(19),
    D => R1IN_3_2F(19),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_156: FDE port map (
    Q => R1IN_3_2F_RETO(20),
    D => R1IN_3_2F(20),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_157: FDE port map (
    Q => R1IN_3_2F_RETO(21),
    D => R1IN_3_2F(21),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_158: FDE port map (
    Q => R1IN_3_2F_RETO(22),
    D => R1IN_3_2F(22),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_159: FDE port map (
    Q => R1IN_3_2F_RETO(23),
    D => R1IN_3_2F(23),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_160: FDE port map (
    Q => R1IN_3_2F_RETO(24),
    D => R1IN_3_2F(24),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_161: FDE port map (
    Q => R1IN_3_2F_RETO(25),
    D => R1IN_3_2F(25),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_162: FDE port map (
    Q => R1IN_3_2F_RETO(26),
    D => R1IN_3_2F(26),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_163: FDE port map (
    Q => R1IN_3_2F_RETO(27),
    D => R1IN_3_2F(27),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_164: FDE port map (
    Q => R1IN_3_2F_RETO(28),
    D => R1IN_3_2F(28),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_165: FDE port map (
    Q => R1IN_3_2F_RETO(29),
    D => R1IN_3_2F(29),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_166: FDE port map (
    Q => R1IN_3_2F_RETO(30),
    D => R1IN_3_2F(30),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_167: FDE port map (
    Q => R1IN_3_2F_RETO(31),
    D => R1IN_3_2F(31),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_168: FDE port map (
    Q => R1IN_3_2F_RETO(32),
    D => R1IN_3_2F(32),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_169: FDE port map (
    Q => R1IN_3_2F_RETO(33),
    D => R1IN_3_2F(33),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_170: FDE port map (
    Q => R1IN_3_2F_RETO(34),
    D => R1IN_3_2F(34),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_171: FDE port map (
    Q => R1IN_3_2F_RETO(35),
    D => R1IN_3_2F(35),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_172: FDE port map (
    Q => R1IN_3_2F_RETO(36),
    D => R1IN_3_2F(36),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_173: FDE port map (
    Q => R1IN_3_2F_RETO(37),
    D => R1IN_3_2F(37),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_174: FDE port map (
    Q => R1IN_3_2F_RETO(38),
    D => R1IN_3_2F(38),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_175: FDE port map (
    Q => R1IN_3_2F_RETO(39),
    D => R1IN_3_2F(39),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_176: FDE port map (
    Q => R1IN_3_2F_RETO(40),
    D => R1IN_3_2F(40),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_177: FDE port map (
    Q => R1IN_3_2F_RETO(41),
    D => R1IN_3_2F(41),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_178: FDE port map (
    Q => R1IN_3_2F_RETO(42),
    D => R1IN_3_2F(42),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_179: FDE port map (
    Q => R1IN_3_2F_RETO(43),
    D => R1IN_3_2F(43),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_91: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO_0(0),
    D => R1IN_4_4_ADD_1F(0),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_92: FDE port map (
    Q => R1IN_4_4_ADD_2_RETO_0,
    D => R1IN_4_4_ADD_2,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_93: FDE port map (
    Q => R1IN_4_4_1F_RETO(18),
    D => R1IN_4_4_1F(18),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_94: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(1),
    D => R1IN_4_4_ADD_1F(1),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_95: FDE port map (
    Q => R1IN_4_4_1F_RETO(19),
    D => R1IN_4_4_1F(19),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_96: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(2),
    D => R1IN_4_4_ADD_1F(2),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_97: FDE port map (
    Q => R1IN_4_4_1F_RETO(20),
    D => R1IN_4_4_1F(20),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_98: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(3),
    D => R1IN_4_4_ADD_1F(3),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_99: FDE port map (
    Q => R1IN_4_4_1F_RETO(21),
    D => R1IN_4_4_1F(21),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_100: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(4),
    D => R1IN_4_4_ADD_1F(4),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_101: FDE port map (
    Q => R1IN_4_4_1F_RETO(22),
    D => R1IN_4_4_1F(22),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_102: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(5),
    D => R1IN_4_4_ADD_1F(5),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_103: FDE port map (
    Q => R1IN_4_4_1F_RETO(23),
    D => R1IN_4_4_1F(23),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_104: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(6),
    D => R1IN_4_4_ADD_1F(6),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_105: FDE port map (
    Q => R1IN_4_4_1F_RETO(24),
    D => R1IN_4_4_1F(24),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_106: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(7),
    D => R1IN_4_4_ADD_1F(7),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_107: FDE port map (
    Q => R1IN_4_4_1F_RETO(25),
    D => R1IN_4_4_1F(25),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_108: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(8),
    D => R1IN_4_4_ADD_1F(8),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_109: FDE port map (
    Q => R1IN_4_4_1F_RETO(26),
    D => R1IN_4_4_1F(26),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_110: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(9),
    D => R1IN_4_4_ADD_1F(9),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_111: FDE port map (
    Q => R1IN_4_4_1F_RETO(27),
    D => R1IN_4_4_1F(27),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_112: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(10),
    D => R1IN_4_4_ADD_1F(10),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_113: FDE port map (
    Q => R1IN_4_4_1F_RETO(28),
    D => R1IN_4_4_1F(28),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_114: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(11),
    D => R1IN_4_4_ADD_1F(11),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_115: FDE port map (
    Q => R1IN_4_4_1F_RETO(29),
    D => R1IN_4_4_1F(29),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_116: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(12),
    D => R1IN_4_4_ADD_1F(12),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_117: FDE port map (
    Q => R1IN_4_4_1F_RETO(30),
    D => R1IN_4_4_1F(30),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_118: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(13),
    D => R1IN_4_4_ADD_1F(13),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_119: FDE port map (
    Q => R1IN_4_4_1F_RETO(31),
    D => R1IN_4_4_1F(31),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_120: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(14),
    D => R1IN_4_4_ADD_1F(14),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_121: FDE port map (
    Q => R1IN_4_4_1F_RETO(32),
    D => R1IN_4_4_1F(32),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_122: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(15),
    D => R1IN_4_4_ADD_1F(15),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_123: FDE port map (
    Q => R1IN_4_4_1F_RETO(33),
    D => R1IN_4_4_1F(33),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_124: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(16),
    D => R1IN_4_4_ADD_1F(16),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_126: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(17),
    D => R1IN_4_4_ADD_1F(17),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_128: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(18),
    D => R1IN_4_4_ADD_1F(18),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_130: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(19),
    D => R1IN_4_4_ADD_1F(19),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_132: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(20),
    D => R1IN_4_4_ADD_1F(20),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_134: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(21),
    D => R1IN_4_4_ADD_1F(21),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_136: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(22),
    D => R1IN_4_4_ADD_1F(22),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_138: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(23),
    D => R1IN_4_4_ADD_1F(23),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_140: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(24),
    D => R1IN_4_4_ADD_1F(24),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_142: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(25),
    D => R1IN_4_4_ADD_1F(25),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_144: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(26),
    D => R1IN_4_4_ADD_1F(26),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_146: FDE port map (
    Q => R1IN_4_4_ADD_1F_RETO(27),
    D => R1IN_4_4_ADD_1F(27),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_60: FDE port map (
    Q => R1IN_2_ADD_1_RETO,
    D => R1IN_2_ADD_1,
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_181: FDE port map (
    Q => R1IN_2_2F_RETO(1),
    D => R1IN_2_2F(1),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_183: FDE port map (
    Q => R1IN_2_2F_RETO(2),
    D => R1IN_2_2F(2),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_185: FDE port map (
    Q => R1IN_2_2F_RETO(3),
    D => R1IN_2_2F(3),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_187: FDE port map (
    Q => R1IN_2_2F_RETO(4),
    D => R1IN_2_2F(4),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_189: FDE port map (
    Q => R1IN_2_2F_RETO(5),
    D => R1IN_2_2F(5),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_191: FDE port map (
    Q => R1IN_2_2F_RETO(6),
    D => R1IN_2_2F(6),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_193: FDE port map (
    Q => R1IN_2_2F_RETO(7),
    D => R1IN_2_2F(7),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_195: FDE port map (
    Q => R1IN_2_2F_RETO(8),
    D => R1IN_2_2F(8),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_197: FDE port map (
    Q => R1IN_2_2F_RETO(9),
    D => R1IN_2_2F(9),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_199: FDE port map (
    Q => R1IN_2_2F_RETO(10),
    D => R1IN_2_2F(10),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_201: FDE port map (
    Q => R1IN_2_2F_RETO(11),
    D => R1IN_2_2F(11),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_203: FDE port map (
    Q => R1IN_2_2F_RETO(12),
    D => R1IN_2_2F(12),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_205: FDE port map (
    Q => R1IN_2_2F_RETO(13),
    D => R1IN_2_2F(13),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_207: FDE port map (
    Q => R1IN_2_2F_RETO(14),
    D => R1IN_2_2F(14),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_209: FDE port map (
    Q => R1IN_2_2F_RETO(15),
    D => R1IN_2_2F(15),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_211: FDE port map (
    Q => R1IN_2_2F_RETO(16),
    D => R1IN_2_2F(16),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_212: FDE port map (
    Q => R1IN_2_2F_RETO(17),
    D => R1IN_2_2F(17),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_213: FDE port map (
    Q => R1IN_2_2F_RETO(18),
    D => R1IN_2_2F(18),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_214: FDE port map (
    Q => R1IN_2_2F_RETO(19),
    D => R1IN_2_2F(19),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_215: FDE port map (
    Q => R1IN_2_2F_RETO(20),
    D => R1IN_2_2F(20),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_216: FDE port map (
    Q => R1IN_2_2F_RETO(21),
    D => R1IN_2_2F(21),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_217: FDE port map (
    Q => R1IN_2_2F_RETO(22),
    D => R1IN_2_2F(22),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_218: FDE port map (
    Q => R1IN_2_2F_RETO(23),
    D => R1IN_2_2F(23),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_219: FDE port map (
    Q => R1IN_2_2F_RETO(24),
    D => R1IN_2_2F(24),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_220: FDE port map (
    Q => R1IN_2_2F_RETO(25),
    D => R1IN_2_2F(25),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_221: FDE port map (
    Q => R1IN_2_2F_RETO(26),
    D => R1IN_2_2F(26),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_222: FDE port map (
    Q => R1IN_2_2F_RETO(27),
    D => R1IN_2_2F(27),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_223: FDE port map (
    Q => R1IN_2_2F_RETO(28),
    D => R1IN_2_2F(28),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_224: FDE port map (
    Q => R1IN_2_2F_RETO(29),
    D => R1IN_2_2F(29),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_225: FDE port map (
    Q => R1IN_2_2F_RETO(30),
    D => R1IN_2_2F(30),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_226: FDE port map (
    Q => R1IN_2_2F_RETO(31),
    D => R1IN_2_2F(31),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_227: FDE port map (
    Q => R1IN_2_2F_RETO(32),
    D => R1IN_2_2F(32),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_228: FDE port map (
    Q => R1IN_2_2F_RETO(33),
    D => R1IN_2_2F(33),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_229: FDE port map (
    Q => R1IN_2_2F_RETO(34),
    D => R1IN_2_2F(34),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_230: FDE port map (
    Q => R1IN_2_2F_RETO(35),
    D => R1IN_2_2F(35),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_231: FDE port map (
    Q => R1IN_2_2F_RETO(36),
    D => R1IN_2_2F(36),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_232: FDE port map (
    Q => R1IN_2_2F_RETO(37),
    D => R1IN_2_2F(37),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_233: FDE port map (
    Q => R1IN_2_2F_RETO(38),
    D => R1IN_2_2F(38),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_234: FDE port map (
    Q => R1IN_2_2F_RETO(39),
    D => R1IN_2_2F(39),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_235: FDE port map (
    Q => R1IN_2_2F_RETO(40),
    D => R1IN_2_2F(40),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_236: FDE port map (
    Q => R1IN_2_2F_RETO(41),
    D => R1IN_2_2F(41),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_237: FDE port map (
    Q => R1IN_2_2F_RETO(42),
    D => R1IN_2_2F(42),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_238: FDE port map (
    Q => R1IN_2_2F_RETO(43),
    D => R1IN_2_2F(43),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_0: FDE port map (
    Q => R1IN_4_3F_RETO(0),
    D => R1IN_4_3F(0),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_62: FDE port map (
    Q => NN_4,
    D => R1IN_4_ADD_1,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_125: FDE port map (
    Q => R1IN_4_2F_RETO(1),
    D => R1IN_4_2F(1),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_127: FDE port map (
    Q => R1IN_4_3F_RETO(1),
    D => R1IN_4_3F(1),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_147: FDE port map (
    Q => R1IN_4_2F_RETO(2),
    D => R1IN_4_2F(2),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_148: FDE port map (
    Q => R1IN_4_3F_RETO(2),
    D => R1IN_4_3F(2),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_149: FDE port map (
    Q => R1IN_4_2F_RETO(3),
    D => R1IN_4_2F(3),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_150: FDE port map (
    Q => R1IN_4_3F_RETO(3),
    D => R1IN_4_3F(3),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_151: FDE port map (
    Q => R1IN_4_2F_RETO(4),
    D => R1IN_4_2F(4),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_152: FDE port map (
    Q => R1IN_4_3F_RETO(4),
    D => R1IN_4_3F(4),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_153: FDE port map (
    Q => R1IN_4_2F_RETO(5),
    D => R1IN_4_2F(5),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_154: FDE port map (
    Q => R1IN_4_3F_RETO(5),
    D => R1IN_4_3F(5),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_155: FDE port map (
    Q => R1IN_4_2F_RETO(6),
    D => R1IN_4_2F(6),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_156: FDE port map (
    Q => R1IN_4_3F_RETO(6),
    D => R1IN_4_3F(6),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_157: FDE port map (
    Q => R1IN_4_2F_RETO(7),
    D => R1IN_4_2F(7),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_158: FDE port map (
    Q => R1IN_4_3F_RETO(7),
    D => R1IN_4_3F(7),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_159: FDE port map (
    Q => R1IN_4_2F_RETO(8),
    D => R1IN_4_2F(8),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_160: FDE port map (
    Q => R1IN_4_3F_RETO(8),
    D => R1IN_4_3F(8),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_161: FDE port map (
    Q => R1IN_4_2F_RETO(9),
    D => R1IN_4_2F(9),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_162: FDE port map (
    Q => R1IN_4_3F_RETO(9),
    D => R1IN_4_3F(9),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_163: FDE port map (
    Q => R1IN_4_2F_RETO(10),
    D => R1IN_4_2F(10),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_164: FDE port map (
    Q => R1IN_4_3F_RETO(10),
    D => R1IN_4_3F(10),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_165: FDE port map (
    Q => R1IN_4_2F_RETO(11),
    D => R1IN_4_2F(11),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_166: FDE port map (
    Q => R1IN_4_3F_RETO(11),
    D => R1IN_4_3F(11),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_167: FDE port map (
    Q => R1IN_4_2F_RETO(12),
    D => R1IN_4_2F(12),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_168: FDE port map (
    Q => R1IN_4_3F_RETO(12),
    D => R1IN_4_3F(12),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_169: FDE port map (
    Q => R1IN_4_2F_RETO(13),
    D => R1IN_4_2F(13),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_170: FDE port map (
    Q => R1IN_4_3F_RETO(13),
    D => R1IN_4_3F(13),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_171: FDE port map (
    Q => R1IN_4_2F_RETO(14),
    D => R1IN_4_2F(14),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_172: FDE port map (
    Q => R1IN_4_3F_RETO(14),
    D => R1IN_4_3F(14),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_173: FDE port map (
    Q => R1IN_4_2F_RETO(15),
    D => R1IN_4_2F(15),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_174: FDE port map (
    Q => R1IN_4_3F_RETO(15),
    D => R1IN_4_3F(15),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_175: FDE port map (
    Q => R1IN_4_2F_RETO(16),
    D => R1IN_4_2F(16),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_176: FDE port map (
    Q => R1IN_4_3F_RETO(16),
    D => R1IN_4_3F(16),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_177: FDE port map (
    Q => R1IN_4_2F_RETO(17),
    D => R1IN_4_2F(17),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_178: FDE port map (
    Q => R1IN_4_3F_RETO(17),
    D => R1IN_4_3F(17),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_179: FDE port map (
    Q => R1IN_4_2F_RETO(18),
    D => R1IN_4_2F(18),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_180: FDE port map (
    Q => R1IN_4_3F_RETO(18),
    D => R1IN_4_3F(18),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_181: FDE port map (
    Q => R1IN_4_2F_RETO(19),
    D => R1IN_4_2F(19),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_182: FDE port map (
    Q => R1IN_4_3F_RETO(19),
    D => R1IN_4_3F(19),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_183: FDE port map (
    Q => R1IN_4_2F_RETO(20),
    D => R1IN_4_2F(20),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_184: FDE port map (
    Q => R1IN_4_3F_RETO(20),
    D => R1IN_4_3F(20),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_185: FDE port map (
    Q => R1IN_4_2F_RETO(21),
    D => R1IN_4_2F(21),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_186: FDE port map (
    Q => R1IN_4_3F_RETO(21),
    D => R1IN_4_3F(21),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_187: FDE port map (
    Q => R1IN_4_2F_RETO(22),
    D => R1IN_4_2F(22),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_188: FDE port map (
    Q => R1IN_4_3F_RETO(22),
    D => R1IN_4_3F(22),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_189: FDE port map (
    Q => R1IN_4_2F_RETO(23),
    D => R1IN_4_2F(23),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_190: FDE port map (
    Q => R1IN_4_3F_RETO(23),
    D => R1IN_4_3F(23),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_191: FDE port map (
    Q => R1IN_4_2F_RETO(24),
    D => R1IN_4_2F(24),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_192: FDE port map (
    Q => R1IN_4_3F_RETO(24),
    D => R1IN_4_3F(24),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_193: FDE port map (
    Q => R1IN_4_2F_RETO(25),
    D => R1IN_4_2F(25),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_194: FDE port map (
    Q => R1IN_4_3F_RETO(25),
    D => R1IN_4_3F(25),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_195: FDE port map (
    Q => R1IN_4_2F_RETO(26),
    D => R1IN_4_2F(26),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_196: FDE port map (
    Q => R1IN_4_3F_RETO(26),
    D => R1IN_4_3F(26),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_197: FDE port map (
    Q => R1IN_4_2F_RETO(27),
    D => R1IN_4_2F(27),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_198: FDE port map (
    Q => R1IN_4_3F_RETO(27),
    D => R1IN_4_3F(27),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_199: FDE port map (
    Q => R1IN_4_2F_RETO(28),
    D => R1IN_4_2F(28),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_200: FDE port map (
    Q => R1IN_4_3F_RETO(28),
    D => R1IN_4_3F(28),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_201: FDE port map (
    Q => R1IN_4_2F_RETO(29),
    D => R1IN_4_2F(29),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_202: FDE port map (
    Q => R1IN_4_3F_RETO(29),
    D => R1IN_4_3F(29),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_203: FDE port map (
    Q => R1IN_4_2F_RETO(30),
    D => R1IN_4_2F(30),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_204: FDE port map (
    Q => R1IN_4_3F_RETO(30),
    D => R1IN_4_3F(30),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_205: FDE port map (
    Q => R1IN_4_2F_RETO(31),
    D => R1IN_4_2F(31),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_206: FDE port map (
    Q => R1IN_4_3F_RETO(31),
    D => R1IN_4_3F(31),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_207: FDE port map (
    Q => R1IN_4_2F_RETO(32),
    D => R1IN_4_2F(32),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_208: FDE port map (
    Q => R1IN_4_3F_RETO(32),
    D => R1IN_4_3F(32),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_209: FDE port map (
    Q => R1IN_4_2F_RETO(33),
    D => R1IN_4_2F(33),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_210: FDE port map (
    Q => R1IN_4_3F_RETO(33),
    D => R1IN_4_3F(33),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_211: FDE port map (
    Q => R1IN_4_2F_RETO(34),
    D => R1IN_4_2F(34),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_212: FDE port map (
    Q => R1IN_4_3F_RETO(34),
    D => R1IN_4_3F(34),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_213: FDE port map (
    Q => R1IN_4_2F_RETO(35),
    D => R1IN_4_2F(35),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_214: FDE port map (
    Q => R1IN_4_3F_RETO(35),
    D => R1IN_4_3F(35),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_215: FDE port map (
    Q => R1IN_4_2F_RETO(36),
    D => R1IN_4_2F(36),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_216: FDE port map (
    Q => R1IN_4_3F_RETO(36),
    D => R1IN_4_3F(36),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_217: FDE port map (
    Q => R1IN_4_2F_RETO(37),
    D => R1IN_4_2F(37),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_218: FDE port map (
    Q => R1IN_4_3F_RETO(37),
    D => R1IN_4_3F(37),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_219: FDE port map (
    Q => R1IN_4_2F_RETO(38),
    D => R1IN_4_2F(38),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_220: FDE port map (
    Q => R1IN_4_3F_RETO(38),
    D => R1IN_4_3F(38),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_221: FDE port map (
    Q => R1IN_4_2F_RETO(39),
    D => R1IN_4_2F(39),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_222: FDE port map (
    Q => R1IN_4_3F_RETO(39),
    D => R1IN_4_3F(39),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_223: FDE port map (
    Q => R1IN_4_2F_RETO(40),
    D => R1IN_4_2F(40),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_224: FDE port map (
    Q => R1IN_4_3F_RETO(40),
    D => R1IN_4_3F(40),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_225: FDE port map (
    Q => R1IN_4_2F_RETO(41),
    D => R1IN_4_2F(41),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_226: FDE port map (
    Q => R1IN_4_3F_RETO(41),
    D => R1IN_4_3F(41),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_227: FDE port map (
    Q => R1IN_4_2F_RETO(42),
    D => R1IN_4_2F(42),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_228: FDE port map (
    Q => R1IN_4_3F_RETO(42),
    D => R1IN_4_3F(42),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_229: FDE port map (
    Q => R1IN_4_2F_RETO(43),
    D => R1IN_4_2F(43),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_230: FDE port map (
    Q => R1IN_4_3F_RETO(43),
    D => R1IN_4_3F(43),
    C => CLK,
    CE => EN);
R1IN_ADD_1_1_CRY_28_Z5102: MUXCY port map (
    DI => R1IN_3(60),
    CI => R1IN_ADD_1_1_CRY_27,
    S => R1IN_ADD_1_1_AXB_28,
    O => R1IN_ADD_1_1_CRY_28);
R1IN_ADD_2_AXB_104_Z5103: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => N_1511,
  I1 => N_1556,
  I2 => R1IN_4_ADD_2_0_CRY_35,
  O => R1IN_ADD_2_AXB_104);
R1IN_4_ADD_1_S_43: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_43,
    CI => R1IN_4_ADD_1_CRY_42,
    O => R1IN_4_ADD_1_RETO(43));
R1IN_4_ADD_1_CRY_43: MUXCY port map (
    DI => R1IN_4_2F_RETO(43),
    CI => R1IN_4_ADD_1_CRY_42,
    S => R1IN_4_ADD_1_AXB_43,
    O => R1IN_4_ADD_1_RETO(44));
R1IN_4_ADD_1_CRY_42_Z5160: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(42),
    CI => R1IN_4_ADD_1_CRY_41,
    S => R1IN_4_ADD_1_AXB_42,
    LO => R1IN_4_ADD_1_CRY_42);
R1IN_4_ADD_1_CRY_41_Z5161: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(41),
    CI => R1IN_4_ADD_1_CRY_40,
    S => R1IN_4_ADD_1_AXB_41,
    LO => R1IN_4_ADD_1_CRY_41);
R1IN_4_ADD_1_S_42: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_42,
    CI => R1IN_4_ADD_1_CRY_41,
    O => R1IN_4_ADD_1_RETO(42));
R1IN_4_ADD_1_CRY_40_Z5163: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(40),
    CI => R1IN_4_ADD_1_CRY_39,
    S => R1IN_4_ADD_1_AXB_40,
    LO => R1IN_4_ADD_1_CRY_40);
R1IN_4_ADD_1_S_41: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_41,
    CI => R1IN_4_ADD_1_CRY_40,
    O => R1IN_4_ADD_1_RETO(41));
R1IN_4_ADD_1_CRY_39_Z5165: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(39),
    CI => R1IN_4_ADD_1_CRY_38,
    S => R1IN_4_ADD_1_AXB_39,
    LO => R1IN_4_ADD_1_CRY_39);
R1IN_4_ADD_1_S_40: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_40,
    CI => R1IN_4_ADD_1_CRY_39,
    O => R1IN_4_ADD_1_RETO(40));
R1IN_4_ADD_1_CRY_38_Z5167: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(38),
    CI => R1IN_4_ADD_1_CRY_37,
    S => R1IN_4_ADD_1_AXB_38,
    LO => R1IN_4_ADD_1_CRY_38);
R1IN_4_ADD_1_S_39: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_39,
    CI => R1IN_4_ADD_1_CRY_38,
    O => R1IN_4_ADD_1_RETO(39));
R1IN_4_ADD_1_CRY_37_Z5169: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(37),
    CI => R1IN_4_ADD_1_CRY_36,
    S => R1IN_4_ADD_1_AXB_37,
    LO => R1IN_4_ADD_1_CRY_37);
R1IN_4_ADD_1_S_38: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_38,
    CI => R1IN_4_ADD_1_CRY_37,
    O => R1IN_4_ADD_1_RETO(38));
R1IN_4_ADD_1_CRY_36_Z5171: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(36),
    CI => R1IN_4_ADD_1_CRY_35,
    S => R1IN_4_ADD_1_AXB_36,
    LO => R1IN_4_ADD_1_CRY_36);
R1IN_4_ADD_1_S_37: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_37,
    CI => R1IN_4_ADD_1_CRY_36,
    O => R1IN_4_ADD_1_RETO(37));
R1IN_4_ADD_1_CRY_35_Z5173: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(35),
    CI => R1IN_4_ADD_1_CRY_34,
    S => R1IN_4_ADD_1_AXB_35,
    LO => R1IN_4_ADD_1_CRY_35);
R1IN_4_ADD_1_S_36: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_36,
    CI => R1IN_4_ADD_1_CRY_35,
    O => R1IN_4_ADD_2_1_RETO);
R1IN_4_ADD_1_CRY_34_Z5175: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(34),
    CI => R1IN_4_ADD_1_CRY_33,
    S => R1IN_4_ADD_1_AXB_34,
    LO => R1IN_4_ADD_1_CRY_34);
R1IN_4_ADD_1_S_35: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_35,
    CI => R1IN_4_ADD_1_CRY_34,
    O => R1IN_4_ADD_1_RETO(35));
R1IN_4_ADD_1_CRY_33_Z5177: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(33),
    CI => R1IN_4_ADD_1_CRY_32,
    S => R1IN_4_ADD_1_AXB_33,
    LO => R1IN_4_ADD_1_CRY_33);
R1IN_4_ADD_1_S_34: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_34,
    CI => R1IN_4_ADD_1_CRY_33,
    O => R1IN_4_ADD_1_RETO(34));
R1IN_4_ADD_1_CRY_32_Z5179: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(32),
    CI => R1IN_4_ADD_1_CRY_31,
    S => R1IN_4_ADD_1_AXB_32,
    LO => R1IN_4_ADD_1_CRY_32);
R1IN_4_ADD_1_S_33: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_33,
    CI => R1IN_4_ADD_1_CRY_32,
    O => R1IN_4_ADD_1_RETO(33));
R1IN_4_ADD_1_CRY_31_Z5181: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(31),
    CI => R1IN_4_ADD_1_CRY_30,
    S => R1IN_4_ADD_1_AXB_31,
    LO => R1IN_4_ADD_1_CRY_31);
R1IN_4_ADD_1_S_32: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_32,
    CI => R1IN_4_ADD_1_CRY_31,
    O => R1IN_4_ADD_1_RETO(32));
R1IN_4_ADD_1_CRY_30_Z5183: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(30),
    CI => R1IN_4_ADD_1_CRY_29,
    S => R1IN_4_ADD_1_AXB_30,
    LO => R1IN_4_ADD_1_CRY_30);
R1IN_4_ADD_1_S_31: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_31,
    CI => R1IN_4_ADD_1_CRY_30,
    O => R1IN_4_ADD_1_RETO(31));
R1IN_4_ADD_1_CRY_29_Z5185: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(29),
    CI => R1IN_4_ADD_1_CRY_28,
    S => R1IN_4_ADD_1_AXB_29,
    LO => R1IN_4_ADD_1_CRY_29);
R1IN_4_ADD_1_S_30: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_30,
    CI => R1IN_4_ADD_1_CRY_29,
    O => R1IN_4_ADD_1_RETO(30));
R1IN_4_ADD_1_CRY_28_Z5187: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(28),
    CI => R1IN_4_ADD_1_CRY_27,
    S => R1IN_4_ADD_1_AXB_28,
    LO => R1IN_4_ADD_1_CRY_28);
R1IN_4_ADD_1_S_29: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_29,
    CI => R1IN_4_ADD_1_CRY_28,
    O => R1IN_4_ADD_1_RETO(29));
R1IN_4_ADD_1_CRY_27_Z5189: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(27),
    CI => R1IN_4_ADD_1_CRY_26,
    S => R1IN_4_ADD_1_AXB_27,
    LO => R1IN_4_ADD_1_CRY_27);
R1IN_4_ADD_1_S_28: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_28,
    CI => R1IN_4_ADD_1_CRY_27,
    O => R1IN_4_ADD_1_RETO(28));
R1IN_4_ADD_1_CRY_26_Z5191: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(26),
    CI => R1IN_4_ADD_1_CRY_25,
    S => R1IN_4_ADD_1_AXB_26,
    LO => R1IN_4_ADD_1_CRY_26);
R1IN_4_ADD_1_S_27: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_27,
    CI => R1IN_4_ADD_1_CRY_26,
    O => R1IN_4_ADD_1_RETO(27));
R1IN_4_ADD_1_CRY_25_Z5193: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(25),
    CI => R1IN_4_ADD_1_CRY_24,
    S => R1IN_4_ADD_1_AXB_25,
    LO => R1IN_4_ADD_1_CRY_25);
R1IN_4_ADD_1_S_26: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_26,
    CI => R1IN_4_ADD_1_CRY_25,
    O => R1IN_4_ADD_1_RETO(26));
R1IN_4_ADD_1_CRY_24_Z5195: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(24),
    CI => R1IN_4_ADD_1_CRY_23,
    S => R1IN_4_ADD_1_AXB_24,
    LO => R1IN_4_ADD_1_CRY_24);
R1IN_4_ADD_1_S_25: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_25,
    CI => R1IN_4_ADD_1_CRY_24,
    O => R1IN_4_ADD_1_RETO(25));
R1IN_4_ADD_1_CRY_23_Z5197: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(23),
    CI => R1IN_4_ADD_1_CRY_22,
    S => R1IN_4_ADD_1_AXB_23,
    LO => R1IN_4_ADD_1_CRY_23);
R1IN_4_ADD_1_S_24: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_24,
    CI => R1IN_4_ADD_1_CRY_23,
    O => R1IN_4_ADD_1_RETO(24));
R1IN_4_ADD_1_CRY_22_Z5199: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(22),
    CI => R1IN_4_ADD_1_CRY_21,
    S => R1IN_4_ADD_1_AXB_22,
    LO => R1IN_4_ADD_1_CRY_22);
R1IN_4_ADD_1_S_23: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_23,
    CI => R1IN_4_ADD_1_CRY_22,
    O => R1IN_4_ADD_1_RETO(23));
R1IN_4_ADD_1_CRY_21_Z5201: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(21),
    CI => R1IN_4_ADD_1_CRY_20,
    S => R1IN_4_ADD_1_AXB_21,
    LO => R1IN_4_ADD_1_CRY_21);
R1IN_4_ADD_1_S_22: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_22,
    CI => R1IN_4_ADD_1_CRY_21,
    O => R1IN_4_ADD_1_RETO(22));
R1IN_4_ADD_1_CRY_20_Z5203: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(20),
    CI => R1IN_4_ADD_1_CRY_19,
    S => R1IN_4_ADD_1_AXB_20,
    LO => R1IN_4_ADD_1_CRY_20);
R1IN_4_ADD_1_S_21: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_21,
    CI => R1IN_4_ADD_1_CRY_20,
    O => R1IN_4_ADD_1_RETO(21));
R1IN_4_ADD_1_CRY_19_Z5205: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(19),
    CI => R1IN_4_ADD_1_CRY_18,
    S => R1IN_4_ADD_1_AXB_19,
    LO => R1IN_4_ADD_1_CRY_19);
R1IN_4_ADD_1_S_20: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_20,
    CI => R1IN_4_ADD_1_CRY_19,
    O => R1IN_4_ADD_1_RETO(20));
R1IN_4_ADD_1_CRY_18_Z5207: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(18),
    CI => R1IN_4_ADD_1_CRY_17,
    S => R1IN_4_ADD_1_AXB_18,
    LO => R1IN_4_ADD_1_CRY_18);
R1IN_4_ADD_1_S_19: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_19,
    CI => R1IN_4_ADD_1_CRY_18,
    O => R1IN_4_ADD_1_RETO(19));
R1IN_4_ADD_1_CRY_17_Z5209: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(17),
    CI => R1IN_4_ADD_1_CRY_16,
    S => R1IN_4_ADD_1_AXB_17,
    LO => R1IN_4_ADD_1_CRY_17);
R1IN_4_ADD_1_S_18: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_18,
    CI => R1IN_4_ADD_1_CRY_17,
    O => R1IN_4_ADD_1_RETO(18));
R1IN_4_ADD_1_CRY_16_Z5211: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(16),
    CI => R1IN_4_ADD_1_CRY_15,
    S => R1IN_4_ADD_1_AXB_16,
    LO => R1IN_4_ADD_1_CRY_16);
R1IN_4_ADD_1_S_17: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_17,
    CI => R1IN_4_ADD_1_CRY_16,
    O => R1IN_4_ADD_1_RETO(17));
R1IN_4_ADD_1_CRY_15_Z5213: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(15),
    CI => R1IN_4_ADD_1_CRY_14,
    S => R1IN_4_ADD_1_AXB_15,
    LO => R1IN_4_ADD_1_CRY_15);
R1IN_4_ADD_1_S_16: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_16,
    CI => R1IN_4_ADD_1_CRY_15,
    O => R1IN_4_ADD_1_RETO(16));
R1IN_4_ADD_1_CRY_14_Z5215: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(14),
    CI => R1IN_4_ADD_1_CRY_13,
    S => R1IN_4_ADD_1_AXB_14,
    LO => R1IN_4_ADD_1_CRY_14);
R1IN_4_ADD_1_S_15: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_15,
    CI => R1IN_4_ADD_1_CRY_14,
    O => R1IN_4_ADD_1_RETO(15));
R1IN_4_ADD_1_CRY_13_Z5217: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(13),
    CI => R1IN_4_ADD_1_CRY_12,
    S => R1IN_4_ADD_1_AXB_13,
    LO => R1IN_4_ADD_1_CRY_13);
R1IN_4_ADD_1_S_14: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_14,
    CI => R1IN_4_ADD_1_CRY_13,
    O => R1IN_4_ADD_1_RETO(14));
R1IN_4_ADD_1_CRY_12_Z5219: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(12),
    CI => R1IN_4_ADD_1_CRY_11,
    S => R1IN_4_ADD_1_AXB_12,
    LO => R1IN_4_ADD_1_CRY_12);
R1IN_4_ADD_1_S_13: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_13,
    CI => R1IN_4_ADD_1_CRY_12,
    O => R1IN_4_ADD_1_RETO(13));
R1IN_4_ADD_1_CRY_11_Z5221: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(11),
    CI => R1IN_4_ADD_1_CRY_10,
    S => R1IN_4_ADD_1_AXB_11,
    LO => R1IN_4_ADD_1_CRY_11);
R1IN_4_ADD_1_S_12: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_12,
    CI => R1IN_4_ADD_1_CRY_11,
    O => R1IN_4_ADD_1_RETO(12));
R1IN_4_ADD_1_CRY_10_Z5223: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(10),
    CI => R1IN_4_ADD_1_CRY_9,
    S => R1IN_4_ADD_1_AXB_10,
    LO => R1IN_4_ADD_1_CRY_10);
R1IN_4_ADD_1_S_11: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_11,
    CI => R1IN_4_ADD_1_CRY_10,
    O => R1IN_4_ADD_1_RETO(11));
R1IN_4_ADD_1_CRY_9_Z5225: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(9),
    CI => R1IN_4_ADD_1_CRY_8,
    S => R1IN_4_ADD_1_AXB_9,
    LO => R1IN_4_ADD_1_CRY_9);
R1IN_4_ADD_1_S_10: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_10,
    CI => R1IN_4_ADD_1_CRY_9,
    O => R1IN_4_ADD_1_RETO(10));
R1IN_4_ADD_1_CRY_8_Z5227: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(8),
    CI => R1IN_4_ADD_1_CRY_7,
    S => R1IN_4_ADD_1_AXB_8,
    LO => R1IN_4_ADD_1_CRY_8);
R1IN_4_ADD_1_S_9: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_9,
    CI => R1IN_4_ADD_1_CRY_8,
    O => R1IN_4_ADD_1_RETO(9));
R1IN_4_ADD_1_CRY_7_Z5229: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(7),
    CI => R1IN_4_ADD_1_CRY_6,
    S => R1IN_4_ADD_1_AXB_7,
    LO => R1IN_4_ADD_1_CRY_7);
R1IN_4_ADD_1_S_8: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_8,
    CI => R1IN_4_ADD_1_CRY_7,
    O => R1IN_4_ADD_1_RETO(8));
R1IN_4_ADD_1_CRY_6_Z5231: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(6),
    CI => R1IN_4_ADD_1_CRY_5,
    S => R1IN_4_ADD_1_AXB_6,
    LO => R1IN_4_ADD_1_CRY_6);
R1IN_4_ADD_1_S_7: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_7,
    CI => R1IN_4_ADD_1_CRY_6,
    O => R1IN_4_ADD_1_RETO(7));
R1IN_4_ADD_1_CRY_5_Z5233: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(5),
    CI => R1IN_4_ADD_1_CRY_4,
    S => R1IN_4_ADD_1_AXB_5,
    LO => R1IN_4_ADD_1_CRY_5);
R1IN_4_ADD_1_S_6: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_6,
    CI => R1IN_4_ADD_1_CRY_5,
    O => R1IN_4_ADD_1_RETO(6));
R1IN_4_ADD_1_CRY_4_Z5235: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(4),
    CI => R1IN_4_ADD_1_CRY_3,
    S => R1IN_4_ADD_1_AXB_4,
    LO => R1IN_4_ADD_1_CRY_4);
R1IN_4_ADD_1_S_5: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_5,
    CI => R1IN_4_ADD_1_CRY_4,
    O => R1IN_4_ADD_1_RETO(5));
R1IN_4_ADD_1_CRY_3_Z5237: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(3),
    CI => R1IN_4_ADD_1_CRY_2,
    S => R1IN_4_ADD_1_AXB_3,
    LO => R1IN_4_ADD_1_CRY_3);
R1IN_4_ADD_1_S_4: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_4,
    CI => R1IN_4_ADD_1_CRY_3,
    O => R1IN_4_ADD_1_RETO(4));
R1IN_4_ADD_1_CRY_2_Z5239: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(2),
    CI => R1IN_4_ADD_1_CRY_1,
    S => R1IN_4_ADD_1_AXB_2,
    LO => R1IN_4_ADD_1_CRY_2);
R1IN_4_ADD_1_S_3: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_3,
    CI => R1IN_4_ADD_1_CRY_2,
    O => R1IN_4_ADD_1_RETO(3));
R1IN_4_ADD_1_CRY_1_Z5241: MUXCY_L port map (
    DI => R1IN_4_2F_RETO(1),
    CI => R1IN_4_ADD_1_CRY_0,
    S => R1IN_4_ADD_1_AXB_1,
    LO => R1IN_4_ADD_1_CRY_1);
R1IN_4_ADD_1_S_2: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_2,
    CI => R1IN_4_ADD_1_CRY_1,
    O => R1IN_4_ADD_1_RETO(2));
R1IN_4_ADD_1_CRY_0_Z5243: MUXCY_L port map (
    DI => NN_4,
    CI => NN_1,
    S => R1IN_4_ADD_2_0_RETO,
    LO => R1IN_4_ADD_1_CRY_0);
R1IN_4_ADD_1_S_1: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_1,
    CI => R1IN_4_ADD_1_CRY_0,
    O => R1IN_4_ADD_1_RETO(1));
R1IN_4_ADD_1_AXB_0: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_3F_RETO(0),
  I1 => NN_4,
  O => R1IN_4_ADD_2_0_RETO);
R1IN_2_ADD_1_S_43: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_43,
    CI => R1IN_2_ADD_1_CRY_42,
    O => R1IN_2_RETO(60));
R1IN_2_ADD_1_AXB_43_Z5320: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F_RETO(43),
  O => R1IN_2_ADD_1_AXB_43);
R1IN_2_ADD_1_CRY_42_Z5321: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_41,
    S => R1IN_2_ADD_1_AXB_42,
    LO => R1IN_2_ADD_1_CRY_42);
R1IN_2_ADD_1_CRY_41_Z5322: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_40,
    S => R1IN_2_ADD_1_AXB_41,
    LO => R1IN_2_ADD_1_CRY_41);
R1IN_2_ADD_1_S_42: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_42,
    CI => R1IN_2_ADD_1_CRY_41,
    O => R1IN_2_RETO(59));
R1IN_2_ADD_1_CRY_40_Z5324: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_39,
    S => R1IN_2_ADD_1_AXB_40,
    LO => R1IN_2_ADD_1_CRY_40);
R1IN_2_ADD_1_S_41: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_41,
    CI => R1IN_2_ADD_1_CRY_40,
    O => R1IN_2_RETO(58));
R1IN_2_ADD_1_CRY_39_Z5326: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_38,
    S => R1IN_2_ADD_1_AXB_39,
    LO => R1IN_2_ADD_1_CRY_39);
R1IN_2_ADD_1_S_40: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_40,
    CI => R1IN_2_ADD_1_CRY_39,
    O => R1IN_2_RETO(57));
R1IN_2_ADD_1_CRY_38_Z5328: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_37,
    S => R1IN_2_ADD_1_AXB_38,
    LO => R1IN_2_ADD_1_CRY_38);
R1IN_2_ADD_1_S_39: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_39,
    CI => R1IN_2_ADD_1_CRY_38,
    O => R1IN_2_RETO(56));
R1IN_2_ADD_1_CRY_37_Z5330: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_36,
    S => R1IN_2_ADD_1_AXB_37,
    LO => R1IN_2_ADD_1_CRY_37);
R1IN_2_ADD_1_S_38: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_38,
    CI => R1IN_2_ADD_1_CRY_37,
    O => R1IN_2_RETO(55));
R1IN_2_ADD_1_CRY_36_Z5332: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_35,
    S => R1IN_2_ADD_1_AXB_36,
    LO => R1IN_2_ADD_1_CRY_36);
R1IN_2_ADD_1_S_37: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_37,
    CI => R1IN_2_ADD_1_CRY_36,
    O => R1IN_2_RETO(54));
R1IN_2_ADD_1_CRY_35_Z5334: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_34,
    S => R1IN_2_ADD_1_AXB_35,
    LO => R1IN_2_ADD_1_CRY_35);
R1IN_2_ADD_1_S_36: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_36,
    CI => R1IN_2_ADD_1_CRY_35,
    O => R1IN_2_RETO(53));
R1IN_2_ADD_1_CRY_34_Z5336: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_33,
    S => R1IN_2_ADD_1_AXB_34,
    LO => R1IN_2_ADD_1_CRY_34);
R1IN_2_ADD_1_S_35: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_35,
    CI => R1IN_2_ADD_1_CRY_34,
    O => R1IN_2_RETO(52));
R1IN_2_ADD_1_CRY_33_Z5338: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_32,
    S => R1IN_2_ADD_1_AXB_33,
    LO => R1IN_2_ADD_1_CRY_33);
R1IN_2_ADD_1_S_34: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_34,
    CI => R1IN_2_ADD_1_CRY_33,
    O => R1IN_2_RETO(51));
R1IN_2_ADD_1_CRY_32_Z5340: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_31,
    S => R1IN_2_ADD_1_AXB_32,
    LO => R1IN_2_ADD_1_CRY_32);
R1IN_2_ADD_1_S_33: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_33,
    CI => R1IN_2_ADD_1_CRY_32,
    O => R1IN_2_RETO(50));
R1IN_2_ADD_1_CRY_31_Z5342: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_30,
    S => R1IN_2_ADD_1_AXB_31,
    LO => R1IN_2_ADD_1_CRY_31);
R1IN_2_ADD_1_S_32: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_32,
    CI => R1IN_2_ADD_1_CRY_31,
    O => R1IN_2_RETO(49));
R1IN_2_ADD_1_CRY_30_Z5344: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_29,
    S => R1IN_2_ADD_1_AXB_30,
    LO => R1IN_2_ADD_1_CRY_30);
R1IN_2_ADD_1_S_31: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_31,
    CI => R1IN_2_ADD_1_CRY_30,
    O => R1IN_2_RETO(48));
R1IN_2_ADD_1_CRY_29_Z5346: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_28,
    S => R1IN_2_ADD_1_AXB_29,
    LO => R1IN_2_ADD_1_CRY_29);
R1IN_2_ADD_1_S_30: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_30,
    CI => R1IN_2_ADD_1_CRY_29,
    O => R1IN_2_RETO(47));
R1IN_2_ADD_1_CRY_28_Z5348: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_27,
    S => R1IN_2_ADD_1_AXB_28,
    LO => R1IN_2_ADD_1_CRY_28);
R1IN_2_ADD_1_S_29: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_29,
    CI => R1IN_2_ADD_1_CRY_28,
    O => R1IN_2_RETO(46));
R1IN_2_ADD_1_CRY_27_Z5350: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_26,
    S => R1IN_2_ADD_1_AXB_27,
    LO => R1IN_2_ADD_1_CRY_27);
R1IN_2_ADD_1_S_28: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_28,
    CI => R1IN_2_ADD_1_CRY_27,
    O => R1IN_2_RETO(45));
R1IN_2_ADD_1_CRY_26_Z5352: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_25,
    S => R1IN_2_ADD_1_AXB_26,
    LO => R1IN_2_ADD_1_CRY_26);
R1IN_2_ADD_1_S_27: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_27,
    CI => R1IN_2_ADD_1_CRY_26,
    O => R1IN_2_RETO(44));
R1IN_2_ADD_1_CRY_25_Z5354: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_24,
    S => R1IN_2_ADD_1_AXB_25,
    LO => R1IN_2_ADD_1_CRY_25);
R1IN_2_ADD_1_S_26: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_26,
    CI => R1IN_2_ADD_1_CRY_25,
    O => R1IN_2_RETO(43));
R1IN_2_ADD_1_CRY_24_Z5356: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_23,
    S => R1IN_2_ADD_1_AXB_24,
    LO => R1IN_2_ADD_1_CRY_24);
R1IN_2_ADD_1_S_25: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_25,
    CI => R1IN_2_ADD_1_CRY_24,
    O => R1IN_2_RETO(42));
R1IN_2_ADD_1_CRY_23_Z5358: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_22,
    S => R1IN_2_ADD_1_AXB_23,
    LO => R1IN_2_ADD_1_CRY_23);
R1IN_2_ADD_1_S_24: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_24,
    CI => R1IN_2_ADD_1_CRY_23,
    O => R1IN_2_RETO(41));
R1IN_2_ADD_1_CRY_22_Z5360: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_21,
    S => R1IN_2_ADD_1_AXB_22,
    LO => R1IN_2_ADD_1_CRY_22);
R1IN_2_ADD_1_S_23: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_23,
    CI => R1IN_2_ADD_1_CRY_22,
    O => R1IN_2_RETO(40));
R1IN_2_ADD_1_CRY_21_Z5362: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_20,
    S => R1IN_2_ADD_1_AXB_21,
    LO => R1IN_2_ADD_1_CRY_21);
R1IN_2_ADD_1_S_22: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_22,
    CI => R1IN_2_ADD_1_CRY_21,
    O => R1IN_2_RETO(39));
R1IN_2_ADD_1_CRY_20_Z5364: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_19,
    S => R1IN_2_ADD_1_AXB_20,
    LO => R1IN_2_ADD_1_CRY_20);
R1IN_2_ADD_1_S_21: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_21,
    CI => R1IN_2_ADD_1_CRY_20,
    O => R1IN_2_RETO(38));
R1IN_2_ADD_1_CRY_19_Z5366: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_18,
    S => R1IN_2_ADD_1_AXB_19,
    LO => R1IN_2_ADD_1_CRY_19);
R1IN_2_ADD_1_S_20: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_20,
    CI => R1IN_2_ADD_1_CRY_19,
    O => R1IN_2_RETO(37));
R1IN_2_ADD_1_CRY_18_Z5368: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_17,
    S => R1IN_2_ADD_1_AXB_18,
    LO => R1IN_2_ADD_1_CRY_18);
R1IN_2_ADD_1_S_19: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_19,
    CI => R1IN_2_ADD_1_CRY_18,
    O => R1IN_2_RETO(36));
R1IN_2_ADD_1_CRY_17_Z5370: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_16,
    S => R1IN_2_ADD_1_AXB_17,
    LO => R1IN_2_ADD_1_CRY_17);
R1IN_2_ADD_1_S_18: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_18,
    CI => R1IN_2_ADD_1_CRY_17,
    O => R1IN_2_RETO(35));
R1IN_2_ADD_1_CRY_16_Z5372: MUXCY_L port map (
    DI => R1IN_2_2F_RETO(16),
    CI => R1IN_2_ADD_1_CRY_15,
    S => R1IN_2_ADD_1_AXB_16,
    LO => R1IN_2_ADD_1_CRY_16);
R1IN_2_ADD_1_S_17: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_17,
    CI => R1IN_2_ADD_1_CRY_16,
    O => R1IN_2_RETO(34));
R1IN_2_ADD_1_CRY_15_Z5374: MUXCY_L port map (
    DI => R1IN_2_2F_RETO(15),
    CI => R1IN_2_ADD_1_CRY_14,
    S => R1IN_2_ADD_1_AXB_15,
    LO => R1IN_2_ADD_1_CRY_15);
R1IN_2_ADD_1_S_16: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_16,
    CI => R1IN_2_ADD_1_CRY_15,
    O => R1IN_2_RETO(33));
R1IN_2_ADD_1_CRY_14_Z5376: MUXCY_L port map (
    DI => R1IN_2_2F_RETO(14),
    CI => R1IN_2_ADD_1_CRY_13,
    S => R1IN_2_ADD_1_AXB_14,
    LO => R1IN_2_ADD_1_CRY_14);
R1IN_2_ADD_1_S_15: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_15,
    CI => R1IN_2_ADD_1_CRY_14,
    O => R1IN_2_RETO(32));
R1IN_2_ADD_1_CRY_13_Z5378: MUXCY_L port map (
    DI => R1IN_2_2F_RETO(13),
    CI => R1IN_2_ADD_1_CRY_12,
    S => R1IN_2_ADD_1_AXB_13,
    LO => R1IN_2_ADD_1_CRY_13);
R1IN_2_ADD_1_S_14: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_14,
    CI => R1IN_2_ADD_1_CRY_13,
    O => R1IN_2_RETO(31));
R1IN_2_ADD_1_CRY_12_Z5380: MUXCY_L port map (
    DI => R1IN_2_2F_RETO(12),
    CI => R1IN_2_ADD_1_CRY_11,
    S => R1IN_2_ADD_1_AXB_12,
    LO => R1IN_2_ADD_1_CRY_12);
R1IN_2_ADD_1_S_13: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_13,
    CI => R1IN_2_ADD_1_CRY_12,
    O => R1IN_2_RETO(30));
R1IN_2_ADD_1_CRY_11_Z5382: MUXCY_L port map (
    DI => R1IN_2_2F_RETO(11),
    CI => R1IN_2_ADD_1_CRY_10,
    S => R1IN_2_ADD_1_AXB_11,
    LO => R1IN_2_ADD_1_CRY_11);
R1IN_2_ADD_1_S_12: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_12,
    CI => R1IN_2_ADD_1_CRY_11,
    O => R1IN_2_RETO(29));
R1IN_2_ADD_1_CRY_10_Z5384: MUXCY_L port map (
    DI => R1IN_2_2F_RETO(10),
    CI => R1IN_2_ADD_1_CRY_9,
    S => R1IN_2_ADD_1_AXB_10,
    LO => R1IN_2_ADD_1_CRY_10);
R1IN_2_ADD_1_S_11: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_11,
    CI => R1IN_2_ADD_1_CRY_10,
    O => R1IN_2_RETO(28));
R1IN_2_ADD_1_CRY_9_Z5386: MUXCY_L port map (
    DI => R1IN_2_2F_RETO(9),
    CI => R1IN_2_ADD_1_CRY_8,
    S => R1IN_2_ADD_1_AXB_9,
    LO => R1IN_2_ADD_1_CRY_9);
R1IN_2_ADD_1_S_10: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_10,
    CI => R1IN_2_ADD_1_CRY_9,
    O => R1IN_2_RETO(27));
R1IN_2_ADD_1_CRY_8_Z5388: MUXCY_L port map (
    DI => R1IN_2_2F_RETO(8),
    CI => R1IN_2_ADD_1_CRY_7,
    S => R1IN_2_ADD_1_AXB_8,
    LO => R1IN_2_ADD_1_CRY_8);
R1IN_2_ADD_1_S_9: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_9,
    CI => R1IN_2_ADD_1_CRY_8,
    O => R1IN_2_RETO(26));
R1IN_2_ADD_1_CRY_7_Z5390: MUXCY_L port map (
    DI => R1IN_2_2F_RETO(7),
    CI => R1IN_2_ADD_1_CRY_6,
    S => R1IN_2_ADD_1_AXB_7,
    LO => R1IN_2_ADD_1_CRY_7);
R1IN_2_ADD_1_S_8: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_8,
    CI => R1IN_2_ADD_1_CRY_7,
    O => R1IN_2_RETO(25));
R1IN_2_ADD_1_CRY_6_Z5392: MUXCY_L port map (
    DI => R1IN_2_2F_RETO(6),
    CI => R1IN_2_ADD_1_CRY_5,
    S => R1IN_2_ADD_1_AXB_6,
    LO => R1IN_2_ADD_1_CRY_6);
R1IN_2_ADD_1_S_7: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_7,
    CI => R1IN_2_ADD_1_CRY_6,
    O => R1IN_2_RETO(24));
R1IN_2_ADD_1_CRY_5_Z5394: MUXCY_L port map (
    DI => R1IN_2_2F_RETO(5),
    CI => R1IN_2_ADD_1_CRY_4,
    S => R1IN_2_ADD_1_AXB_5,
    LO => R1IN_2_ADD_1_CRY_5);
R1IN_2_ADD_1_S_6: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_6,
    CI => R1IN_2_ADD_1_CRY_5,
    O => R1IN_2_RETO(23));
R1IN_2_ADD_1_CRY_4_Z5396: MUXCY_L port map (
    DI => R1IN_2_2F_RETO(4),
    CI => R1IN_2_ADD_1_CRY_3,
    S => R1IN_2_ADD_1_AXB_4,
    LO => R1IN_2_ADD_1_CRY_4);
R1IN_2_ADD_1_S_5: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_5,
    CI => R1IN_2_ADD_1_CRY_4,
    O => R1IN_2_RETO(22));
R1IN_2_ADD_1_CRY_3_Z5398: MUXCY_L port map (
    DI => R1IN_2_2F_RETO(3),
    CI => R1IN_2_ADD_1_CRY_2,
    S => R1IN_2_ADD_1_AXB_3,
    LO => R1IN_2_ADD_1_CRY_3);
R1IN_2_ADD_1_S_4: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_4,
    CI => R1IN_2_ADD_1_CRY_3,
    O => R1IN_2_RETO(21));
R1IN_2_ADD_1_CRY_2_Z5400: MUXCY_L port map (
    DI => R1IN_2_2F_RETO(2),
    CI => R1IN_2_ADD_1_CRY_1,
    S => R1IN_2_ADD_1_AXB_2,
    LO => R1IN_2_ADD_1_CRY_2);
R1IN_2_ADD_1_S_3: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_3,
    CI => R1IN_2_ADD_1_CRY_2,
    O => R1IN_2_RETO(20));
R1IN_2_ADD_1_CRY_1_Z5402: MUXCY_L port map (
    DI => R1IN_2_2F_RETO(1),
    CI => R1IN_2_ADD_1_CRY_0,
    S => R1IN_2_ADD_1_AXB_1,
    LO => R1IN_2_ADD_1_CRY_1);
R1IN_2_ADD_1_S_2: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_2,
    CI => R1IN_2_ADD_1_CRY_1,
    O => R1IN_2_RETO(19));
R1IN_2_ADD_1_CRY_0_Z5404: MUXCY_L port map (
    DI => R1IN_2_ADD_1_RETO,
    CI => NN_1,
    S => R1IN_2_RETO(17),
    LO => R1IN_2_ADD_1_CRY_0);
R1IN_2_ADD_1_S_1: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_1,
    CI => R1IN_2_ADD_1_CRY_0,
    O => R1IN_2_RETO(18));
R1IN_2_ADD_1_AXB_0: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F_RETO(17),
  I1 => R1IN_2_ADD_1_RETO,
  O => R1IN_2_RETO(17));
R1IN_4_ADD_2_0_AXB_1_Z5879: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F_RETO(18),
  I1 => R1IN_4_ADD_1_RETO(1),
  LO => R1IN_4_ADD_2_0_AXB_1);
R1IN_4_ADD_2_0_AXB_2_Z5880: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F_RETO(19),
  I1 => R1IN_4_ADD_1_RETO(2),
  LO => R1IN_4_ADD_2_0_AXB_2);
R1IN_4_ADD_2_0_AXB_3_Z5881: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F_RETO(20),
  I1 => R1IN_4_ADD_1_RETO(3),
  LO => R1IN_4_ADD_2_0_AXB_3);
R1IN_4_ADD_2_0_AXB_4_Z5882: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F_RETO(21),
  I1 => R1IN_4_ADD_1_RETO(4),
  LO => R1IN_4_ADD_2_0_AXB_4);
R1IN_4_ADD_2_0_AXB_5_Z5883: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F_RETO(22),
  I1 => R1IN_4_ADD_1_RETO(5),
  LO => R1IN_4_ADD_2_0_AXB_5);
R1IN_4_ADD_2_0_AXB_6_Z5884: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F_RETO(23),
  I1 => R1IN_4_ADD_1_RETO(6),
  LO => R1IN_4_ADD_2_0_AXB_6);
R1IN_4_ADD_2_0_AXB_7_Z5885: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F_RETO(24),
  I1 => R1IN_4_ADD_1_RETO(7),
  LO => R1IN_4_ADD_2_0_AXB_7);
R1IN_4_ADD_2_0_AXB_8_Z5886: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F_RETO(25),
  I1 => R1IN_4_ADD_1_RETO(8),
  LO => R1IN_4_ADD_2_0_AXB_8);
R1IN_4_ADD_2_0_AXB_9_Z5887: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F_RETO(26),
  I1 => R1IN_4_ADD_1_RETO(9),
  LO => R1IN_4_ADD_2_0_AXB_9);
R1IN_4_ADD_2_0_AXB_10_Z5888: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F_RETO(27),
  I1 => R1IN_4_ADD_1_RETO(10),
  LO => R1IN_4_ADD_2_0_AXB_10);
R1IN_4_ADD_2_0_AXB_11_Z5889: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F_RETO(28),
  I1 => R1IN_4_ADD_1_RETO(11),
  LO => R1IN_4_ADD_2_0_AXB_11);
R1IN_4_ADD_2_0_AXB_12_Z5890: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F_RETO(29),
  I1 => R1IN_4_ADD_1_RETO(12),
  LO => R1IN_4_ADD_2_0_AXB_12);
R1IN_4_ADD_2_0_AXB_13_Z5891: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F_RETO(30),
  I1 => R1IN_4_ADD_1_RETO(13),
  LO => R1IN_4_ADD_2_0_AXB_13);
R1IN_4_ADD_2_0_AXB_14_Z5892: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F_RETO(31),
  I1 => R1IN_4_ADD_1_RETO(14),
  LO => R1IN_4_ADD_2_0_AXB_14);
R1IN_4_ADD_2_0_AXB_15_Z5893: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F_RETO(32),
  I1 => R1IN_4_ADD_1_RETO(15),
  LO => R1IN_4_ADD_2_0_AXB_15);
R1IN_4_ADD_2_0_AXB_16_Z5894: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F_RETO(33),
  I1 => R1IN_4_ADD_1_RETO(16),
  LO => R1IN_4_ADD_2_0_AXB_16);
R1IN_4_ADD_2_0_AXB_17_Z5895: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F_RETO(0),
  I1 => R1IN_4_ADD_1_RETO(17),
  LO => R1IN_4_ADD_2_0_AXB_17);
R1IN_4_ADD_2_0_AXB_18_Z5896: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F_RETO(1),
  I1 => R1IN_4_ADD_1_RETO(18),
  LO => R1IN_4_ADD_2_0_AXB_18);
R1IN_4_ADD_2_0_AXB_19_Z5897: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F_RETO(2),
  I1 => R1IN_4_ADD_1_RETO(19),
  LO => R1IN_4_ADD_2_0_AXB_19);
R1IN_4_ADD_2_0_AXB_20_Z5898: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F_RETO(3),
  I1 => R1IN_4_ADD_1_RETO(20),
  LO => R1IN_4_ADD_2_0_AXB_20);
R1IN_4_ADD_2_0_AXB_21_Z5899: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F_RETO(4),
  I1 => R1IN_4_ADD_1_RETO(21),
  LO => R1IN_4_ADD_2_0_AXB_21);
R1IN_4_ADD_2_0_AXB_22_Z5900: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F_RETO(5),
  I1 => R1IN_4_ADD_1_RETO(22),
  LO => R1IN_4_ADD_2_0_AXB_22);
R1IN_4_ADD_2_0_AXB_23_Z5901: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F_RETO(6),
  I1 => R1IN_4_ADD_1_RETO(23),
  LO => R1IN_4_ADD_2_0_AXB_23);
R1IN_4_ADD_2_0_AXB_24_Z5902: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F_RETO(7),
  I1 => R1IN_4_ADD_1_RETO(24),
  LO => R1IN_4_ADD_2_0_AXB_24);
R1IN_4_ADD_2_0_AXB_25_Z5903: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F_RETO(8),
  I1 => R1IN_4_ADD_1_RETO(25),
  LO => R1IN_4_ADD_2_0_AXB_25);
R1IN_4_ADD_2_0_AXB_26_Z5904: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F_RETO(9),
  I1 => R1IN_4_ADD_1_RETO(26),
  LO => R1IN_4_ADD_2_0_AXB_26);
R1IN_4_ADD_2_0_AXB_27_Z5905: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F_RETO(10),
  I1 => R1IN_4_ADD_1_RETO(27),
  LO => R1IN_4_ADD_2_0_AXB_27);
R1IN_4_ADD_2_0_AXB_28_Z5906: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F_RETO(11),
  I1 => R1IN_4_ADD_1_RETO(28),
  LO => R1IN_4_ADD_2_0_AXB_28);
R1IN_4_ADD_2_0_AXB_29_Z5907: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F_RETO(12),
  I1 => R1IN_4_ADD_1_RETO(29),
  LO => R1IN_4_ADD_2_0_AXB_29);
R1IN_4_ADD_2_0_AXB_30_Z5908: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F_RETO(13),
  I1 => R1IN_4_ADD_1_RETO(30),
  LO => R1IN_4_ADD_2_0_AXB_30);
R1IN_4_ADD_2_0_AXB_31_Z5909: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F_RETO(14),
  I1 => R1IN_4_ADD_1_RETO(31),
  LO => R1IN_4_ADD_2_0_AXB_31);
R1IN_4_ADD_2_0_AXB_32_Z5910: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F_RETO(15),
  I1 => R1IN_4_ADD_1_RETO(32),
  LO => R1IN_4_ADD_2_0_AXB_32);
R1IN_4_ADD_2_0_AXB_33_Z5911: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F_RETO(16),
  I1 => R1IN_4_ADD_1_RETO(33),
  LO => R1IN_4_ADD_2_0_AXB_33);
R1IN_4_ADD_2_0_AXB_34_Z5912: LUT3_L 
generic map(
  INIT => X"96"
)
port map (
  I0 => R1IN_4_4_ADD_1F_RETO(0),
  I1 => R1IN_4_4_ADD_2_RETO,
  I2 => R1IN_4_ADD_1_RETO(34),
  LO => R1IN_4_ADD_2_0_AXB_34);
R1IN_4_ADD_2_0_AXB_35_Z5913: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(18),
  I1 => R1IN_4_ADD_1_RETO(35),
  LO => R1IN_4_ADD_2_0_AXB_35);
R1IN_ADD_1_0_AXB_1_Z5914: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F_RETO(1),
  I1 => R1IN_3F_RETO(1),
  LO => R1IN_ADD_1_0_AXB_1);
R1IN_ADD_1_0_AXB_2_Z5915: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F_RETO(2),
  I1 => R1IN_3F_RETO(2),
  LO => R1IN_ADD_1_0_AXB_2);
R1IN_ADD_1_0_AXB_3_Z5916: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F_RETO(3),
  I1 => R1IN_3F_RETO(3),
  LO => R1IN_ADD_1_0_AXB_3);
R1IN_ADD_1_0_AXB_4_Z5917: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F_RETO(4),
  I1 => R1IN_3F_RETO(4),
  LO => R1IN_ADD_1_0_AXB_4);
R1IN_ADD_1_0_AXB_5_Z5918: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F_RETO(5),
  I1 => R1IN_3F_RETO(5),
  LO => R1IN_ADD_1_0_AXB_5);
R1IN_ADD_1_0_AXB_6_Z5919: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F_RETO(6),
  I1 => R1IN_3F_RETO(6),
  LO => R1IN_ADD_1_0_AXB_6);
R1IN_ADD_1_0_AXB_7_Z5920: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F_RETO(7),
  I1 => R1IN_3F_RETO(7),
  LO => R1IN_ADD_1_0_AXB_7);
R1IN_ADD_1_0_AXB_8_Z5921: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F_RETO(8),
  I1 => R1IN_3F_RETO(8),
  LO => R1IN_ADD_1_0_AXB_8);
R1IN_ADD_1_0_AXB_9_Z5922: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F_RETO(9),
  I1 => R1IN_3F_RETO(9),
  LO => R1IN_ADD_1_0_AXB_9);
R1IN_ADD_1_0_AXB_10_Z5923: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F_RETO(10),
  I1 => R1IN_3F_RETO(10),
  LO => R1IN_ADD_1_0_AXB_10);
R1IN_ADD_1_0_AXB_11_Z5924: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F_RETO(11),
  I1 => R1IN_3F_RETO(11),
  LO => R1IN_ADD_1_0_AXB_11);
R1IN_ADD_1_0_AXB_12_Z5925: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F_RETO(12),
  I1 => R1IN_3F_RETO(12),
  LO => R1IN_ADD_1_0_AXB_12);
R1IN_ADD_1_0_AXB_13_Z5926: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F_RETO(13),
  I1 => R1IN_3F_RETO(13),
  LO => R1IN_ADD_1_0_AXB_13);
R1IN_ADD_1_0_AXB_14_Z5927: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F_RETO(14),
  I1 => R1IN_3F_RETO(14),
  LO => R1IN_ADD_1_0_AXB_14);
R1IN_ADD_1_0_AXB_15_Z5928: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F_RETO(15),
  I1 => R1IN_3F_RETO(15),
  LO => R1IN_ADD_1_0_AXB_15);
R1IN_ADD_1_0_AXB_16_Z5929: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F_RETO(16),
  I1 => R1IN_3F_RETO(16),
  LO => R1IN_ADD_1_0_AXB_16);
R1IN_ADD_1_0_AXB_17_Z5930: LUT3_L 
generic map(
  INIT => X"96"
)
port map (
  I0 => R1IN_2_RETO(17),
  I1 => R1IN_3_1F_RETO(17),
  I2 => R1IN_3_ADD_1_RETO,
  LO => R1IN_ADD_1_0_AXB_17);
R1IN_ADD_1_0_AXB_18_Z5931: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(18),
  I1 => R1IN_3(18),
  LO => R1IN_ADD_1_0_AXB_18);
R1IN_ADD_1_0_AXB_19_Z5932: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(19),
  I1 => R1IN_3(19),
  LO => R1IN_ADD_1_0_AXB_19);
R1IN_ADD_1_0_AXB_20_Z5933: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(20),
  I1 => R1IN_3(20),
  LO => R1IN_ADD_1_0_AXB_20);
R1IN_ADD_1_0_AXB_21_Z5934: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(21),
  I1 => R1IN_3(21),
  LO => R1IN_ADD_1_0_AXB_21);
R1IN_ADD_1_0_AXB_22_Z5935: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(22),
  I1 => R1IN_3(22),
  LO => R1IN_ADD_1_0_AXB_22);
R1IN_ADD_1_0_AXB_23_Z5936: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(23),
  I1 => R1IN_3(23),
  LO => R1IN_ADD_1_0_AXB_23);
R1IN_ADD_1_0_AXB_24_Z5937: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(24),
  I1 => R1IN_3(24),
  LO => R1IN_ADD_1_0_AXB_24);
R1IN_ADD_1_0_AXB_25_Z5938: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(25),
  I1 => R1IN_3(25),
  LO => R1IN_ADD_1_0_AXB_25);
R1IN_ADD_1_0_AXB_26_Z5939: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(26),
  I1 => R1IN_3(26),
  LO => R1IN_ADD_1_0_AXB_26);
R1IN_ADD_1_0_AXB_27_Z5940: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(27),
  I1 => R1IN_3(27),
  LO => R1IN_ADD_1_0_AXB_27);
R1IN_ADD_1_0_AXB_28_Z5941: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(28),
  I1 => R1IN_3(28),
  LO => R1IN_ADD_1_0_AXB_28);
R1IN_ADD_1_0_AXB_29_Z5942: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(29),
  I1 => R1IN_3(29),
  LO => R1IN_ADD_1_0_AXB_29);
R1IN_ADD_1_0_AXB_30_Z5943: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(30),
  I1 => R1IN_3(30),
  LO => R1IN_ADD_1_0_AXB_30);
R1IN_ADD_1_0_AXB_31_Z5944: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(31),
  I1 => R1IN_3(31),
  LO => R1IN_ADD_1_0_AXB_31);
R1IN_ADD_2_AXB_0: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_ADD_1(0),
  I1 => R1IN_ADD_2,
  O => NN_3);
R1IN_4_4_ADD_2_AXB_36_Z5946: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4_4F_RETO(19),
  O => R1IN_4_4_ADD_2_AXB_36);
R1IN_3_ADD_1_AXB_43_Z5947: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F_RETO(43),
  O => R1IN_3_ADD_1_AXB_43);
R1IN_3_ADD_1_AXB_0: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F_RETO_0(17),
  I1 => R1IN_3_ADD_1_RETO_0,
  O => R1IN_3(17));
R1IN_ADD_1_1_0_AXB_0_Z5949: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(32),
  I1 => R1IN_3(32),
  O => R1IN_ADD_1_1_0_AXB_0);
R1IN_ADD_1_1_AXB_0_Z5950: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_RETO(32),
  I1 => R1IN_3(32),
  O => R1IN_ADD_1_1_AXB_0);
R1IN_ADD_1_0_AXB_0: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F_RETO(0),
  I1 => R1IN_3F_RETO(0),
  O => R1IN_ADD_1(0));
R1IN_4_ADD_2_1_0_AXB_34_Z5952: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(53),
  O => R1IN_4_ADD_2_1_0_AXB_34);
R1IN_4_ADD_2_1_0_AXB_0_Z5953: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(19),
  I1 => R1IN_4_ADD_2_1_RETO,
  O => R1IN_4_ADD_2_1_0_AXB_0);
R1IN_4_ADD_2_1_AXB_34_Z5954: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(53),
  O => R1IN_4_ADD_2_1_AXB_34);
R1IN_4_ADD_2_1_AXB_0_Z5955: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(19),
  I1 => R1IN_4_ADD_2_1_RETO,
  O => R1IN_4_ADD_2_1_AXB_0);
R1IN_4_ADD_2_0_AXB_0: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F_RETO(17),
  I1 => R1IN_4_ADD_2_0_RETO,
  O => R1IN_4(17));
R1IN_ADD_2_S_104: XORCY port map (
    LI => R1IN_ADD_2_AXB_104,
    CI => R1IN_ADD_2_CRY_103,
    O => PRODUCT(121));
R1IN_ADD_2_S_103: XORCY port map (
    LI => R1IN_ADD_2_AXB_103,
    CI => R1IN_ADD_2_CRY_102,
    O => PRODUCT(120));
R1IN_ADD_2_CRY_103_Z5959: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_102,
    S => R1IN_ADD_2_AXB_103,
    LO => R1IN_ADD_2_CRY_103);
R1IN_ADD_2_S_102: XORCY port map (
    LI => R1IN_ADD_2_AXB_102,
    CI => R1IN_ADD_2_CRY_101,
    O => PRODUCT(119));
R1IN_ADD_2_CRY_102_Z5961: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_101,
    S => R1IN_ADD_2_AXB_102,
    LO => R1IN_ADD_2_CRY_102);
R1IN_ADD_2_S_101: XORCY port map (
    LI => R1IN_ADD_2_AXB_101,
    CI => R1IN_ADD_2_CRY_100,
    O => PRODUCT(118));
R1IN_ADD_2_CRY_101_Z5963: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_100,
    S => R1IN_ADD_2_AXB_101,
    LO => R1IN_ADD_2_CRY_101);
R1IN_ADD_2_S_100: XORCY port map (
    LI => R1IN_ADD_2_AXB_100,
    CI => R1IN_ADD_2_CRY_99,
    O => PRODUCT(117));
R1IN_ADD_2_CRY_100_Z5965: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_99,
    S => R1IN_ADD_2_AXB_100,
    LO => R1IN_ADD_2_CRY_100);
R1IN_ADD_2_S_99: XORCY port map (
    LI => R1IN_ADD_2_AXB_99,
    CI => R1IN_ADD_2_CRY_98,
    O => PRODUCT(116));
R1IN_ADD_2_CRY_99_Z5967: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_98,
    S => R1IN_ADD_2_AXB_99,
    LO => R1IN_ADD_2_CRY_99);
R1IN_ADD_2_S_98: XORCY port map (
    LI => R1IN_ADD_2_AXB_98,
    CI => R1IN_ADD_2_CRY_97,
    O => PRODUCT(115));
R1IN_ADD_2_CRY_98_Z5969: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_97,
    S => R1IN_ADD_2_AXB_98,
    LO => R1IN_ADD_2_CRY_98);
R1IN_ADD_2_S_97: XORCY port map (
    LI => R1IN_ADD_2_AXB_97,
    CI => R1IN_ADD_2_CRY_96,
    O => PRODUCT(114));
R1IN_ADD_2_CRY_97_Z5971: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_96,
    S => R1IN_ADD_2_AXB_97,
    LO => R1IN_ADD_2_CRY_97);
R1IN_ADD_2_S_96: XORCY port map (
    LI => R1IN_ADD_2_AXB_96,
    CI => R1IN_ADD_2_CRY_95,
    O => PRODUCT(113));
R1IN_ADD_2_CRY_96_Z5973: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_95,
    S => R1IN_ADD_2_AXB_96,
    LO => R1IN_ADD_2_CRY_96);
R1IN_ADD_2_S_95: XORCY port map (
    LI => R1IN_ADD_2_AXB_95,
    CI => R1IN_ADD_2_CRY_94,
    O => PRODUCT(112));
R1IN_ADD_2_CRY_95_Z5975: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_94,
    S => R1IN_ADD_2_AXB_95,
    LO => R1IN_ADD_2_CRY_95);
R1IN_ADD_2_S_94: XORCY port map (
    LI => R1IN_ADD_2_AXB_94,
    CI => R1IN_ADD_2_CRY_93,
    O => PRODUCT(111));
R1IN_ADD_2_CRY_94_Z5977: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_93,
    S => R1IN_ADD_2_AXB_94,
    LO => R1IN_ADD_2_CRY_94);
R1IN_ADD_2_S_93: XORCY port map (
    LI => R1IN_ADD_2_AXB_93,
    CI => R1IN_ADD_2_CRY_92,
    O => PRODUCT(110));
R1IN_ADD_2_CRY_93_Z5979: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_92,
    S => R1IN_ADD_2_AXB_93,
    LO => R1IN_ADD_2_CRY_93);
R1IN_ADD_2_S_92: XORCY port map (
    LI => R1IN_ADD_2_AXB_92,
    CI => R1IN_ADD_2_CRY_91,
    O => PRODUCT(109));
R1IN_ADD_2_CRY_92_Z5981: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_91,
    S => R1IN_ADD_2_AXB_92,
    LO => R1IN_ADD_2_CRY_92);
R1IN_ADD_2_S_91: XORCY port map (
    LI => R1IN_ADD_2_AXB_91,
    CI => R1IN_ADD_2_CRY_90,
    O => PRODUCT(108));
R1IN_ADD_2_CRY_91_Z5983: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_90,
    S => R1IN_ADD_2_AXB_91,
    LO => R1IN_ADD_2_CRY_91);
R1IN_ADD_2_S_90: XORCY port map (
    LI => R1IN_ADD_2_AXB_90,
    CI => R1IN_ADD_2_CRY_89,
    O => PRODUCT(107));
R1IN_ADD_2_CRY_90_Z5985: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_89,
    S => R1IN_ADD_2_AXB_90,
    LO => R1IN_ADD_2_CRY_90);
R1IN_ADD_2_S_89: XORCY port map (
    LI => R1IN_ADD_2_AXB_89,
    CI => R1IN_ADD_2_CRY_88,
    O => PRODUCT(106));
R1IN_ADD_2_CRY_89_Z5987: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_88,
    S => R1IN_ADD_2_AXB_89,
    LO => R1IN_ADD_2_CRY_89);
R1IN_ADD_2_S_88: XORCY port map (
    LI => R1IN_ADD_2_AXB_88,
    CI => R1IN_ADD_2_CRY_87,
    O => PRODUCT(105));
R1IN_ADD_2_CRY_88_Z5989: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_87,
    S => R1IN_ADD_2_AXB_88,
    LO => R1IN_ADD_2_CRY_88);
R1IN_ADD_2_S_87: XORCY port map (
    LI => R1IN_ADD_2_AXB_87,
    CI => R1IN_ADD_2_CRY_86,
    O => PRODUCT(104));
R1IN_ADD_2_CRY_87_Z5991: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_86,
    S => R1IN_ADD_2_AXB_87,
    LO => R1IN_ADD_2_CRY_87);
R1IN_ADD_2_S_86: XORCY port map (
    LI => R1IN_ADD_2_AXB_86,
    CI => R1IN_ADD_2_CRY_85,
    O => PRODUCT(103));
R1IN_ADD_2_CRY_86_Z5993: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_85,
    S => R1IN_ADD_2_AXB_86,
    LO => R1IN_ADD_2_CRY_86);
R1IN_ADD_2_S_85: XORCY port map (
    LI => R1IN_ADD_2_AXB_85,
    CI => R1IN_ADD_2_CRY_84,
    O => PRODUCT(102));
R1IN_ADD_2_CRY_85_Z5995: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_84,
    S => R1IN_ADD_2_AXB_85,
    LO => R1IN_ADD_2_CRY_85);
R1IN_ADD_2_S_84: XORCY port map (
    LI => R1IN_ADD_2_AXB_84,
    CI => R1IN_ADD_2_CRY_83,
    O => PRODUCT(101));
R1IN_ADD_2_CRY_84_Z5997: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_83,
    S => R1IN_ADD_2_AXB_84,
    LO => R1IN_ADD_2_CRY_84);
R1IN_ADD_2_S_83: XORCY port map (
    LI => R1IN_ADD_2_AXB_83,
    CI => R1IN_ADD_2_CRY_82,
    O => PRODUCT(100));
R1IN_ADD_2_CRY_83_Z5999: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_82,
    S => R1IN_ADD_2_AXB_83,
    LO => R1IN_ADD_2_CRY_83);
R1IN_ADD_2_S_82: XORCY port map (
    LI => R1IN_ADD_2_AXB_82,
    CI => R1IN_ADD_2_CRY_81,
    O => PRODUCT(99));
R1IN_ADD_2_CRY_82_Z6001: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_81,
    S => R1IN_ADD_2_AXB_82,
    LO => R1IN_ADD_2_CRY_82);
R1IN_ADD_2_S_81: XORCY port map (
    LI => R1IN_ADD_2_AXB_81,
    CI => R1IN_ADD_2_CRY_80,
    O => PRODUCT(98));
R1IN_ADD_2_CRY_81_Z6003: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_80,
    S => R1IN_ADD_2_AXB_81,
    LO => R1IN_ADD_2_CRY_81);
R1IN_ADD_2_S_80: XORCY port map (
    LI => R1IN_ADD_2_AXB_80,
    CI => R1IN_ADD_2_CRY_79,
    O => PRODUCT(97));
R1IN_ADD_2_CRY_80_Z6005: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_79,
    S => R1IN_ADD_2_AXB_80,
    LO => R1IN_ADD_2_CRY_80);
R1IN_ADD_2_S_79: XORCY port map (
    LI => R1IN_ADD_2_AXB_79,
    CI => R1IN_ADD_2_CRY_78,
    O => PRODUCT(96));
R1IN_ADD_2_CRY_79_Z6007: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_78,
    S => R1IN_ADD_2_AXB_79,
    LO => R1IN_ADD_2_CRY_79);
R1IN_ADD_2_S_78: XORCY port map (
    LI => R1IN_ADD_2_AXB_78,
    CI => R1IN_ADD_2_CRY_77,
    O => PRODUCT(95));
R1IN_ADD_2_CRY_78_Z6009: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_77,
    S => R1IN_ADD_2_AXB_78,
    LO => R1IN_ADD_2_CRY_78);
R1IN_ADD_2_S_77: XORCY port map (
    LI => R1IN_ADD_2_AXB_77,
    CI => R1IN_ADD_2_CRY_76,
    O => PRODUCT(94));
R1IN_ADD_2_CRY_77_Z6011: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_76,
    S => R1IN_ADD_2_AXB_77,
    LO => R1IN_ADD_2_CRY_77);
R1IN_ADD_2_S_76: XORCY port map (
    LI => R1IN_ADD_2_AXB_76,
    CI => R1IN_ADD_2_CRY_75,
    O => PRODUCT(93));
R1IN_ADD_2_CRY_76_Z6013: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_75,
    S => R1IN_ADD_2_AXB_76,
    LO => R1IN_ADD_2_CRY_76);
R1IN_ADD_2_S_75: XORCY port map (
    LI => R1IN_ADD_2_AXB_75,
    CI => R1IN_ADD_2_CRY_74,
    O => PRODUCT(92));
R1IN_ADD_2_CRY_75_Z6015: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_74,
    S => R1IN_ADD_2_AXB_75,
    LO => R1IN_ADD_2_CRY_75);
R1IN_ADD_2_S_74: XORCY port map (
    LI => R1IN_ADD_2_AXB_74,
    CI => R1IN_ADD_2_CRY_73,
    O => PRODUCT(91));
R1IN_ADD_2_CRY_74_Z6017: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_73,
    S => R1IN_ADD_2_AXB_74,
    LO => R1IN_ADD_2_CRY_74);
R1IN_ADD_2_S_73: XORCY port map (
    LI => R1IN_ADD_2_AXB_73,
    CI => R1IN_ADD_2_CRY_72,
    O => PRODUCT(90));
R1IN_ADD_2_CRY_73_Z6019: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_72,
    S => R1IN_ADD_2_AXB_73,
    LO => R1IN_ADD_2_CRY_73);
R1IN_ADD_2_S_72: XORCY port map (
    LI => R1IN_ADD_2_AXB_72,
    CI => R1IN_ADD_2_CRY_71,
    O => PRODUCT(89));
R1IN_ADD_2_CRY_72_Z6021: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_71,
    S => R1IN_ADD_2_AXB_72,
    LO => R1IN_ADD_2_CRY_72);
R1IN_ADD_2_S_71: XORCY port map (
    LI => R1IN_ADD_2_AXB_71,
    CI => R1IN_ADD_2_CRY_70,
    O => PRODUCT(88));
R1IN_ADD_2_CRY_71_Z6023: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_70,
    S => R1IN_ADD_2_AXB_71,
    LO => R1IN_ADD_2_CRY_71);
R1IN_ADD_2_S_70: XORCY port map (
    LI => R1IN_ADD_2_AXB_70,
    CI => R1IN_ADD_2_CRY_69,
    O => PRODUCT(87));
R1IN_ADD_2_CRY_70_Z6025: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_69,
    S => R1IN_ADD_2_AXB_70,
    LO => R1IN_ADD_2_CRY_70);
R1IN_ADD_2_S_69: XORCY port map (
    LI => R1IN_ADD_2_AXB_69,
    CI => R1IN_ADD_2_CRY_68,
    O => PRODUCT(86));
R1IN_ADD_2_CRY_69_Z6027: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_68,
    S => R1IN_ADD_2_AXB_69,
    LO => R1IN_ADD_2_CRY_69);
R1IN_ADD_2_S_68: XORCY port map (
    LI => R1IN_ADD_2_AXB_68,
    CI => R1IN_ADD_2_CRY_67,
    O => PRODUCT(85));
R1IN_ADD_2_CRY_68_Z6029: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_67,
    S => R1IN_ADD_2_AXB_68,
    LO => R1IN_ADD_2_CRY_68);
R1IN_ADD_2_S_67: XORCY port map (
    LI => R1IN_ADD_2_AXB_67,
    CI => R1IN_ADD_2_CRY_66,
    O => PRODUCT(84));
R1IN_ADD_2_CRY_67_Z6031: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_66,
    S => R1IN_ADD_2_AXB_67,
    LO => R1IN_ADD_2_CRY_67);
R1IN_ADD_2_S_66: XORCY port map (
    LI => R1IN_ADD_2_AXB_66,
    CI => R1IN_ADD_2_CRY_65,
    O => PRODUCT(83));
R1IN_ADD_2_CRY_66_Z6033: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_65,
    S => R1IN_ADD_2_AXB_66,
    LO => R1IN_ADD_2_CRY_66);
R1IN_ADD_2_S_65: XORCY port map (
    LI => R1IN_ADD_2_AXB_65,
    CI => R1IN_ADD_2_CRY_64,
    O => PRODUCT(82));
R1IN_ADD_2_CRY_65_Z6035: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_64,
    S => R1IN_ADD_2_AXB_65,
    LO => R1IN_ADD_2_CRY_65);
R1IN_ADD_2_S_64: XORCY port map (
    LI => R1IN_ADD_2_AXB_64,
    CI => R1IN_ADD_2_CRY_63,
    O => PRODUCT(81));
R1IN_ADD_2_CRY_64_Z6037: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_63,
    S => R1IN_ADD_2_AXB_64,
    LO => R1IN_ADD_2_CRY_64);
R1IN_ADD_2_S_63: XORCY port map (
    LI => R1IN_ADD_2_AXB_63,
    CI => R1IN_ADD_2_CRY_62,
    O => PRODUCT(80));
R1IN_ADD_2_CRY_63_Z6039: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_62,
    S => R1IN_ADD_2_AXB_63,
    LO => R1IN_ADD_2_CRY_63);
R1IN_ADD_2_S_62: XORCY port map (
    LI => R1IN_ADD_2_AXB_62,
    CI => R1IN_ADD_2_CRY_61,
    O => PRODUCT(79));
R1IN_ADD_2_CRY_62_Z6041: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_CRY_61,
    S => R1IN_ADD_2_AXB_62,
    LO => R1IN_ADD_2_CRY_62);
R1IN_ADD_2_S_61: XORCY port map (
    LI => R1IN_ADD_2_AXB_61,
    CI => R1IN_ADD_2_CRY_60,
    O => PRODUCT(78));
R1IN_ADD_2_CRY_61_Z6043: MUXCY_L port map (
    DI => R1IN_4(44),
    CI => R1IN_ADD_2_CRY_60,
    S => R1IN_ADD_2_AXB_61,
    LO => R1IN_ADD_2_CRY_61);
R1IN_ADD_2_S_60: XORCY port map (
    LI => R1IN_ADD_2_AXB_60,
    CI => R1IN_ADD_2_CRY_59,
    O => PRODUCT(77));
R1IN_ADD_2_CRY_60_Z6045: MUXCY_L port map (
    DI => R1IN_4(43),
    CI => R1IN_ADD_2_CRY_59,
    S => R1IN_ADD_2_AXB_60,
    LO => R1IN_ADD_2_CRY_60);
R1IN_ADD_2_S_59: XORCY port map (
    LI => R1IN_ADD_2_AXB_59,
    CI => R1IN_ADD_2_CRY_58,
    O => PRODUCT(76));
R1IN_ADD_2_CRY_59_Z6047: MUXCY_L port map (
    DI => R1IN_4(42),
    CI => R1IN_ADD_2_CRY_58,
    S => R1IN_ADD_2_AXB_59,
    LO => R1IN_ADD_2_CRY_59);
R1IN_ADD_2_S_58: XORCY port map (
    LI => R1IN_ADD_2_AXB_58,
    CI => R1IN_ADD_2_CRY_57,
    O => PRODUCT(75));
R1IN_ADD_2_CRY_58_Z6049: MUXCY_L port map (
    DI => R1IN_4(41),
    CI => R1IN_ADD_2_CRY_57,
    S => R1IN_ADD_2_AXB_58,
    LO => R1IN_ADD_2_CRY_58);
R1IN_ADD_2_S_57: XORCY port map (
    LI => R1IN_ADD_2_AXB_57,
    CI => R1IN_ADD_2_CRY_56,
    O => PRODUCT(74));
R1IN_ADD_2_CRY_57_Z6051: MUXCY_L port map (
    DI => R1IN_4(40),
    CI => R1IN_ADD_2_CRY_56,
    S => R1IN_ADD_2_AXB_57,
    LO => R1IN_ADD_2_CRY_57);
R1IN_ADD_2_S_56: XORCY port map (
    LI => R1IN_ADD_2_AXB_56,
    CI => R1IN_ADD_2_CRY_55,
    O => PRODUCT(73));
R1IN_ADD_2_CRY_56_Z6053: MUXCY_L port map (
    DI => R1IN_4(39),
    CI => R1IN_ADD_2_CRY_55,
    S => R1IN_ADD_2_AXB_56,
    LO => R1IN_ADD_2_CRY_56);
R1IN_ADD_2_S_55: XORCY port map (
    LI => R1IN_ADD_2_AXB_55,
    CI => R1IN_ADD_2_CRY_54,
    O => PRODUCT(72));
R1IN_ADD_2_CRY_55_Z6055: MUXCY_L port map (
    DI => R1IN_4(38),
    CI => R1IN_ADD_2_CRY_54,
    S => R1IN_ADD_2_AXB_55,
    LO => R1IN_ADD_2_CRY_55);
R1IN_ADD_2_S_54: XORCY port map (
    LI => R1IN_ADD_2_AXB_54,
    CI => R1IN_ADD_2_CRY_53,
    O => PRODUCT(71));
R1IN_ADD_2_CRY_54_Z6057: MUXCY_L port map (
    DI => R1IN_4(37),
    CI => R1IN_ADD_2_CRY_53,
    S => R1IN_ADD_2_AXB_54,
    LO => R1IN_ADD_2_CRY_54);
R1IN_ADD_2_S_53: XORCY port map (
    LI => R1IN_ADD_2_AXB_53,
    CI => R1IN_ADD_2_CRY_52,
    O => PRODUCT(70));
R1IN_ADD_2_CRY_53_Z6059: MUXCY_L port map (
    DI => R1IN_4(36),
    CI => R1IN_ADD_2_CRY_52,
    S => R1IN_ADD_2_AXB_53,
    LO => R1IN_ADD_2_CRY_53);
R1IN_ADD_2_S_52: XORCY port map (
    LI => R1IN_ADD_2_AXB_52,
    CI => R1IN_ADD_2_CRY_51,
    O => PRODUCT(69));
R1IN_ADD_2_CRY_52_Z6061: MUXCY_L port map (
    DI => R1IN_4(35),
    CI => R1IN_ADD_2_CRY_51,
    S => R1IN_ADD_2_AXB_52,
    LO => R1IN_ADD_2_CRY_52);
R1IN_ADD_2_S_51: XORCY port map (
    LI => R1IN_ADD_2_AXB_51,
    CI => R1IN_ADD_2_CRY_50,
    O => PRODUCT(68));
R1IN_ADD_2_CRY_51_Z6063: MUXCY_L port map (
    DI => R1IN_4(34),
    CI => R1IN_ADD_2_CRY_50,
    S => R1IN_ADD_2_AXB_51,
    LO => R1IN_ADD_2_CRY_51);
R1IN_ADD_2_S_50: XORCY port map (
    LI => R1IN_ADD_2_AXB_50,
    CI => R1IN_ADD_2_CRY_49,
    O => PRODUCT(67));
R1IN_ADD_2_CRY_50_Z6065: MUXCY_L port map (
    DI => R1IN_4(33),
    CI => R1IN_ADD_2_CRY_49,
    S => R1IN_ADD_2_AXB_50,
    LO => R1IN_ADD_2_CRY_50);
R1IN_ADD_2_S_49: XORCY port map (
    LI => R1IN_ADD_2_AXB_49,
    CI => R1IN_ADD_2_CRY_48,
    O => PRODUCT(66));
R1IN_ADD_2_CRY_49_Z6067: MUXCY_L port map (
    DI => R1IN_4(32),
    CI => R1IN_ADD_2_CRY_48,
    S => R1IN_ADD_2_AXB_49,
    LO => R1IN_ADD_2_CRY_49);
R1IN_ADD_2_S_48: XORCY port map (
    LI => R1IN_ADD_2_AXB_48,
    CI => R1IN_ADD_2_CRY_47,
    O => PRODUCT(65));
R1IN_ADD_2_CRY_48_Z6069: MUXCY_L port map (
    DI => R1IN_4(31),
    CI => R1IN_ADD_2_CRY_47,
    S => R1IN_ADD_2_AXB_48,
    LO => R1IN_ADD_2_CRY_48);
R1IN_ADD_2_S_47: XORCY port map (
    LI => R1IN_ADD_2_AXB_47,
    CI => R1IN_ADD_2_CRY_46,
    O => PRODUCT(64));
R1IN_ADD_2_CRY_47_Z6071: MUXCY_L port map (
    DI => R1IN_4(30),
    CI => R1IN_ADD_2_CRY_46,
    S => R1IN_ADD_2_AXB_47,
    LO => R1IN_ADD_2_CRY_47);
R1IN_ADD_2_S_46: XORCY port map (
    LI => R1IN_ADD_2_AXB_46,
    CI => R1IN_ADD_2_CRY_45,
    O => PRODUCT(63));
R1IN_ADD_2_CRY_46_Z6073: MUXCY_L port map (
    DI => R1IN_4(29),
    CI => R1IN_ADD_2_CRY_45,
    S => R1IN_ADD_2_AXB_46,
    LO => R1IN_ADD_2_CRY_46);
R1IN_ADD_2_S_45: XORCY port map (
    LI => R1IN_ADD_2_AXB_45,
    CI => R1IN_ADD_2_CRY_44,
    O => PRODUCT(62));
R1IN_ADD_2_CRY_45_Z6075: MUXCY_L port map (
    DI => R1IN_4(28),
    CI => R1IN_ADD_2_CRY_44,
    S => R1IN_ADD_2_AXB_45,
    LO => R1IN_ADD_2_CRY_45);
R1IN_ADD_2_S_44: XORCY port map (
    LI => R1IN_ADD_2_AXB_44,
    CI => R1IN_ADD_2_CRY_43,
    O => PRODUCT(61));
R1IN_ADD_2_CRY_44_Z6077: MUXCY_L port map (
    DI => R1IN_4(27),
    CI => R1IN_ADD_2_CRY_43,
    S => R1IN_ADD_2_AXB_44,
    LO => R1IN_ADD_2_CRY_44);
R1IN_ADD_2_S_43: XORCY port map (
    LI => R1IN_ADD_2_AXB_43,
    CI => R1IN_ADD_2_CRY_42,
    O => PRODUCT(60));
R1IN_ADD_2_CRY_43_Z6079: MUXCY_L port map (
    DI => R1IN_4(26),
    CI => R1IN_ADD_2_CRY_42,
    S => R1IN_ADD_2_AXB_43,
    LO => R1IN_ADD_2_CRY_43);
R1IN_ADD_2_S_42: XORCY port map (
    LI => R1IN_ADD_2_AXB_42,
    CI => R1IN_ADD_2_CRY_41,
    O => PRODUCT(59));
R1IN_ADD_2_CRY_42_Z6081: MUXCY_L port map (
    DI => R1IN_4(25),
    CI => R1IN_ADD_2_CRY_41,
    S => R1IN_ADD_2_AXB_42,
    LO => R1IN_ADD_2_CRY_42);
R1IN_ADD_2_S_41: XORCY port map (
    LI => R1IN_ADD_2_AXB_41,
    CI => R1IN_ADD_2_CRY_40,
    O => PRODUCT(58));
R1IN_ADD_2_CRY_41_Z6083: MUXCY_L port map (
    DI => R1IN_4(24),
    CI => R1IN_ADD_2_CRY_40,
    S => R1IN_ADD_2_AXB_41,
    LO => R1IN_ADD_2_CRY_41);
R1IN_ADD_2_S_40: XORCY port map (
    LI => R1IN_ADD_2_AXB_40,
    CI => R1IN_ADD_2_CRY_39,
    O => PRODUCT(57));
R1IN_ADD_2_CRY_40_Z6085: MUXCY_L port map (
    DI => R1IN_4(23),
    CI => R1IN_ADD_2_CRY_39,
    S => R1IN_ADD_2_AXB_40,
    LO => R1IN_ADD_2_CRY_40);
R1IN_ADD_2_S_39: XORCY port map (
    LI => R1IN_ADD_2_AXB_39,
    CI => R1IN_ADD_2_CRY_38,
    O => PRODUCT(56));
R1IN_ADD_2_CRY_39_Z6087: MUXCY_L port map (
    DI => R1IN_4(22),
    CI => R1IN_ADD_2_CRY_38,
    S => R1IN_ADD_2_AXB_39,
    LO => R1IN_ADD_2_CRY_39);
R1IN_ADD_2_S_38: XORCY port map (
    LI => R1IN_ADD_2_AXB_38,
    CI => R1IN_ADD_2_CRY_37,
    O => PRODUCT(55));
R1IN_ADD_2_CRY_38_Z6089: MUXCY_L port map (
    DI => R1IN_4(21),
    CI => R1IN_ADD_2_CRY_37,
    S => R1IN_ADD_2_AXB_38,
    LO => R1IN_ADD_2_CRY_38);
R1IN_ADD_2_S_37: XORCY port map (
    LI => R1IN_ADD_2_AXB_37,
    CI => R1IN_ADD_2_CRY_36,
    O => PRODUCT(54));
R1IN_ADD_2_CRY_37_Z6091: MUXCY_L port map (
    DI => R1IN_4(20),
    CI => R1IN_ADD_2_CRY_36,
    S => R1IN_ADD_2_AXB_37,
    LO => R1IN_ADD_2_CRY_37);
R1IN_ADD_2_S_36: XORCY port map (
    LI => R1IN_ADD_2_AXB_36,
    CI => R1IN_ADD_2_CRY_35,
    O => PRODUCT(53));
R1IN_ADD_2_CRY_36_Z6093: MUXCY_L port map (
    DI => R1IN_4(19),
    CI => R1IN_ADD_2_CRY_35,
    S => R1IN_ADD_2_AXB_36,
    LO => R1IN_ADD_2_CRY_36);
R1IN_ADD_2_S_35: XORCY port map (
    LI => R1IN_ADD_2_AXB_35,
    CI => R1IN_ADD_2_CRY_34,
    O => PRODUCT(52));
R1IN_ADD_2_CRY_35_Z6095: MUXCY_L port map (
    DI => R1IN_4(18),
    CI => R1IN_ADD_2_CRY_34,
    S => R1IN_ADD_2_AXB_35,
    LO => R1IN_ADD_2_CRY_35);
R1IN_ADD_2_S_34: XORCY port map (
    LI => R1IN_ADD_2_AXB_34,
    CI => R1IN_ADD_2_CRY_33,
    O => PRODUCT(51));
R1IN_ADD_2_CRY_34_Z6097: MUXCY_L port map (
    DI => R1IN_4(17),
    CI => R1IN_ADD_2_CRY_33,
    S => R1IN_ADD_2_AXB_34,
    LO => R1IN_ADD_2_CRY_34);
R1IN_ADD_2_S_33: XORCY port map (
    LI => R1IN_ADD_2_AXB_33,
    CI => R1IN_ADD_2_CRY_32,
    O => PRODUCT(50));
R1IN_ADD_2_CRY_33_Z6099: MUXCY_L port map (
    DI => R1IN_4FF(16),
    CI => R1IN_ADD_2_CRY_32,
    S => R1IN_ADD_2_AXB_33,
    LO => R1IN_ADD_2_CRY_33);
R1IN_ADD_2_S_32: XORCY port map (
    LI => R1IN_ADD_2_AXB_32,
    CI => R1IN_ADD_2_CRY_31,
    O => PRODUCT(49));
R1IN_ADD_2_CRY_32_Z6101: MUXCY_L port map (
    DI => R1IN_4FF(15),
    CI => R1IN_ADD_2_CRY_31,
    S => R1IN_ADD_2_AXB_32,
    LO => R1IN_ADD_2_CRY_32);
R1IN_ADD_2_S_31: XORCY port map (
    LI => R1IN_ADD_2_AXB_31,
    CI => R1IN_ADD_2_CRY_30,
    O => PRODUCT(48));
R1IN_ADD_2_CRY_31_Z6103: MUXCY_L port map (
    DI => R1IN_4FF(14),
    CI => R1IN_ADD_2_CRY_30,
    S => R1IN_ADD_2_AXB_31,
    LO => R1IN_ADD_2_CRY_31);
R1IN_ADD_2_S_30: XORCY port map (
    LI => R1IN_ADD_2_AXB_30,
    CI => R1IN_ADD_2_CRY_29,
    O => PRODUCT(47));
R1IN_ADD_2_CRY_30_Z6105: MUXCY_L port map (
    DI => R1IN_4FF(13),
    CI => R1IN_ADD_2_CRY_29,
    S => R1IN_ADD_2_AXB_30,
    LO => R1IN_ADD_2_CRY_30);
R1IN_ADD_2_S_29: XORCY port map (
    LI => R1IN_ADD_2_AXB_29,
    CI => R1IN_ADD_2_CRY_28,
    O => PRODUCT(46));
R1IN_ADD_2_CRY_29_Z6107: MUXCY_L port map (
    DI => R1IN_4FF(12),
    CI => R1IN_ADD_2_CRY_28,
    S => R1IN_ADD_2_AXB_29,
    LO => R1IN_ADD_2_CRY_29);
R1IN_ADD_2_S_28: XORCY port map (
    LI => R1IN_ADD_2_AXB_28,
    CI => R1IN_ADD_2_CRY_27,
    O => PRODUCT(45));
R1IN_ADD_2_CRY_28_Z6109: MUXCY_L port map (
    DI => R1IN_4FF(11),
    CI => R1IN_ADD_2_CRY_27,
    S => R1IN_ADD_2_AXB_28,
    LO => R1IN_ADD_2_CRY_28);
R1IN_ADD_2_S_27: XORCY port map (
    LI => R1IN_ADD_2_AXB_27,
    CI => R1IN_ADD_2_CRY_26,
    O => PRODUCT(44));
R1IN_ADD_2_CRY_27_Z6111: MUXCY_L port map (
    DI => R1IN_4FF(10),
    CI => R1IN_ADD_2_CRY_26,
    S => R1IN_ADD_2_AXB_27,
    LO => R1IN_ADD_2_CRY_27);
R1IN_ADD_2_S_26: XORCY port map (
    LI => R1IN_ADD_2_AXB_26,
    CI => R1IN_ADD_2_CRY_25,
    O => PRODUCT(43));
R1IN_ADD_2_CRY_26_Z6113: MUXCY_L port map (
    DI => R1IN_4FF(9),
    CI => R1IN_ADD_2_CRY_25,
    S => R1IN_ADD_2_AXB_26,
    LO => R1IN_ADD_2_CRY_26);
R1IN_ADD_2_S_25: XORCY port map (
    LI => R1IN_ADD_2_AXB_25,
    CI => R1IN_ADD_2_CRY_24,
    O => PRODUCT(42));
R1IN_ADD_2_CRY_25_Z6115: MUXCY_L port map (
    DI => R1IN_4FF(8),
    CI => R1IN_ADD_2_CRY_24,
    S => R1IN_ADD_2_AXB_25,
    LO => R1IN_ADD_2_CRY_25);
R1IN_ADD_2_S_24: XORCY port map (
    LI => R1IN_ADD_2_AXB_24,
    CI => R1IN_ADD_2_CRY_23,
    O => PRODUCT(41));
R1IN_ADD_2_CRY_24_Z6117: MUXCY_L port map (
    DI => R1IN_4FF(7),
    CI => R1IN_ADD_2_CRY_23,
    S => R1IN_ADD_2_AXB_24,
    LO => R1IN_ADD_2_CRY_24);
R1IN_ADD_2_S_23: XORCY port map (
    LI => R1IN_ADD_2_AXB_23,
    CI => R1IN_ADD_2_CRY_22,
    O => PRODUCT(40));
R1IN_ADD_2_CRY_23_Z6119: MUXCY_L port map (
    DI => R1IN_4FF(6),
    CI => R1IN_ADD_2_CRY_22,
    S => R1IN_ADD_2_AXB_23,
    LO => R1IN_ADD_2_CRY_23);
R1IN_ADD_2_S_22: XORCY port map (
    LI => R1IN_ADD_2_AXB_22,
    CI => R1IN_ADD_2_CRY_21,
    O => PRODUCT(39));
R1IN_ADD_2_CRY_22_Z6121: MUXCY_L port map (
    DI => R1IN_4FF(5),
    CI => R1IN_ADD_2_CRY_21,
    S => R1IN_ADD_2_AXB_22,
    LO => R1IN_ADD_2_CRY_22);
R1IN_ADD_2_S_21: XORCY port map (
    LI => R1IN_ADD_2_AXB_21,
    CI => R1IN_ADD_2_CRY_20,
    O => PRODUCT(38));
R1IN_ADD_2_CRY_21_Z6123: MUXCY_L port map (
    DI => R1IN_4FF(4),
    CI => R1IN_ADD_2_CRY_20,
    S => R1IN_ADD_2_AXB_21,
    LO => R1IN_ADD_2_CRY_21);
R1IN_ADD_2_S_20: XORCY port map (
    LI => R1IN_ADD_2_AXB_20,
    CI => R1IN_ADD_2_CRY_19,
    O => PRODUCT(37));
R1IN_ADD_2_CRY_20_Z6125: MUXCY_L port map (
    DI => R1IN_4FF(3),
    CI => R1IN_ADD_2_CRY_19,
    S => R1IN_ADD_2_AXB_20,
    LO => R1IN_ADD_2_CRY_20);
R1IN_ADD_2_S_19: XORCY port map (
    LI => R1IN_ADD_2_AXB_19,
    CI => R1IN_ADD_2_CRY_18,
    O => PRODUCT(36));
R1IN_ADD_2_CRY_19_Z6127: MUXCY_L port map (
    DI => R1IN_4FF(2),
    CI => R1IN_ADD_2_CRY_18,
    S => R1IN_ADD_2_AXB_19,
    LO => R1IN_ADD_2_CRY_19);
R1IN_ADD_2_S_18: XORCY port map (
    LI => R1IN_ADD_2_AXB_18,
    CI => R1IN_ADD_2_CRY_17,
    O => PRODUCT(35));
R1IN_ADD_2_CRY_18_Z6129: MUXCY_L port map (
    DI => R1IN_4FF(1),
    CI => R1IN_ADD_2_CRY_17,
    S => R1IN_ADD_2_AXB_18,
    LO => R1IN_ADD_2_CRY_18);
R1IN_ADD_2_S_17: XORCY port map (
    LI => R1IN_ADD_2_AXB_17,
    CI => R1IN_ADD_2_CRY_16,
    O => PRODUCT(34));
R1IN_ADD_2_CRY_17_Z6131: MUXCY_L port map (
    DI => R1IN_4FF(0),
    CI => R1IN_ADD_2_CRY_16,
    S => R1IN_ADD_2_AXB_17,
    LO => R1IN_ADD_2_CRY_17);
R1IN_ADD_2_S_16: XORCY port map (
    LI => R1IN_ADD_2_AXB_16,
    CI => R1IN_ADD_2_CRY_15,
    O => PRODUCT(33));
R1IN_ADD_2_CRY_16_Z6133: MUXCY_L port map (
    DI => R1IN_1FF(33),
    CI => R1IN_ADD_2_CRY_15,
    S => R1IN_ADD_2_AXB_16,
    LO => R1IN_ADD_2_CRY_16);
R1IN_ADD_2_S_15: XORCY port map (
    LI => R1IN_ADD_2_AXB_15,
    CI => R1IN_ADD_2_CRY_14,
    O => PRODUCT(32));
R1IN_ADD_2_CRY_15_Z6135: MUXCY_L port map (
    DI => R1IN_1FF(32),
    CI => R1IN_ADD_2_CRY_14,
    S => R1IN_ADD_2_AXB_15,
    LO => R1IN_ADD_2_CRY_15);
R1IN_ADD_2_S_14: XORCY port map (
    LI => R1IN_ADD_2_AXB_14,
    CI => R1IN_ADD_2_CRY_13,
    O => PRODUCT(31));
R1IN_ADD_2_CRY_14_Z6137: MUXCY_L port map (
    DI => R1IN_1FF(31),
    CI => R1IN_ADD_2_CRY_13,
    S => R1IN_ADD_2_AXB_14,
    LO => R1IN_ADD_2_CRY_14);
R1IN_ADD_2_S_13: XORCY port map (
    LI => R1IN_ADD_2_AXB_13,
    CI => R1IN_ADD_2_CRY_12,
    O => PRODUCT(30));
R1IN_ADD_2_CRY_13_Z6139: MUXCY_L port map (
    DI => R1IN_1FF(30),
    CI => R1IN_ADD_2_CRY_12,
    S => R1IN_ADD_2_AXB_13,
    LO => R1IN_ADD_2_CRY_13);
R1IN_ADD_2_S_12: XORCY port map (
    LI => R1IN_ADD_2_AXB_12,
    CI => R1IN_ADD_2_CRY_11,
    O => PRODUCT(29));
R1IN_ADD_2_CRY_12_Z6141: MUXCY_L port map (
    DI => R1IN_1FF(29),
    CI => R1IN_ADD_2_CRY_11,
    S => R1IN_ADD_2_AXB_12,
    LO => R1IN_ADD_2_CRY_12);
R1IN_ADD_2_S_11: XORCY port map (
    LI => R1IN_ADD_2_AXB_11,
    CI => R1IN_ADD_2_CRY_10,
    O => PRODUCT(28));
R1IN_ADD_2_CRY_11_Z6143: MUXCY_L port map (
    DI => R1IN_1FF(28),
    CI => R1IN_ADD_2_CRY_10,
    S => R1IN_ADD_2_AXB_11,
    LO => R1IN_ADD_2_CRY_11);
R1IN_ADD_2_S_10: XORCY port map (
    LI => R1IN_ADD_2_AXB_10,
    CI => R1IN_ADD_2_CRY_9,
    O => PRODUCT(27));
R1IN_ADD_2_CRY_10_Z6145: MUXCY_L port map (
    DI => R1IN_1FF(27),
    CI => R1IN_ADD_2_CRY_9,
    S => R1IN_ADD_2_AXB_10,
    LO => R1IN_ADD_2_CRY_10);
R1IN_ADD_2_S_9: XORCY port map (
    LI => R1IN_ADD_2_AXB_9,
    CI => R1IN_ADD_2_CRY_8,
    O => PRODUCT(26));
R1IN_ADD_2_CRY_9_Z6147: MUXCY_L port map (
    DI => R1IN_1FF(26),
    CI => R1IN_ADD_2_CRY_8,
    S => R1IN_ADD_2_AXB_9,
    LO => R1IN_ADD_2_CRY_9);
R1IN_ADD_2_S_8: XORCY port map (
    LI => R1IN_ADD_2_AXB_8,
    CI => R1IN_ADD_2_CRY_7,
    O => PRODUCT(25));
R1IN_ADD_2_CRY_8_Z6149: MUXCY_L port map (
    DI => R1IN_1FF(25),
    CI => R1IN_ADD_2_CRY_7,
    S => R1IN_ADD_2_AXB_8,
    LO => R1IN_ADD_2_CRY_8);
R1IN_ADD_2_S_7: XORCY port map (
    LI => R1IN_ADD_2_AXB_7,
    CI => R1IN_ADD_2_CRY_6,
    O => PRODUCT(24));
R1IN_ADD_2_CRY_7_Z6151: MUXCY_L port map (
    DI => R1IN_1FF(24),
    CI => R1IN_ADD_2_CRY_6,
    S => R1IN_ADD_2_AXB_7,
    LO => R1IN_ADD_2_CRY_7);
R1IN_ADD_2_S_6: XORCY port map (
    LI => R1IN_ADD_2_AXB_6,
    CI => R1IN_ADD_2_CRY_5,
    O => PRODUCT(23));
R1IN_ADD_2_CRY_6_Z6153: MUXCY_L port map (
    DI => R1IN_1FF(23),
    CI => R1IN_ADD_2_CRY_5,
    S => R1IN_ADD_2_AXB_6,
    LO => R1IN_ADD_2_CRY_6);
R1IN_ADD_2_S_5: XORCY port map (
    LI => R1IN_ADD_2_AXB_5,
    CI => R1IN_ADD_2_CRY_4,
    O => PRODUCT(22));
R1IN_ADD_2_CRY_5_Z6155: MUXCY_L port map (
    DI => R1IN_1FF(22),
    CI => R1IN_ADD_2_CRY_4,
    S => R1IN_ADD_2_AXB_5,
    LO => R1IN_ADD_2_CRY_5);
R1IN_ADD_2_S_4: XORCY port map (
    LI => R1IN_ADD_2_AXB_4,
    CI => R1IN_ADD_2_CRY_3,
    O => PRODUCT(21));
R1IN_ADD_2_CRY_4_Z6157: MUXCY_L port map (
    DI => R1IN_1FF(21),
    CI => R1IN_ADD_2_CRY_3,
    S => R1IN_ADD_2_AXB_4,
    LO => R1IN_ADD_2_CRY_4);
R1IN_ADD_2_S_3: XORCY port map (
    LI => R1IN_ADD_2_AXB_3,
    CI => R1IN_ADD_2_CRY_2,
    O => PRODUCT(20));
R1IN_ADD_2_CRY_3_Z6159: MUXCY_L port map (
    DI => R1IN_1FF(20),
    CI => R1IN_ADD_2_CRY_2,
    S => R1IN_ADD_2_AXB_3,
    LO => R1IN_ADD_2_CRY_3);
R1IN_ADD_2_S_2: XORCY port map (
    LI => R1IN_ADD_2_AXB_2,
    CI => R1IN_ADD_2_CRY_1,
    O => PRODUCT(19));
R1IN_ADD_2_CRY_2_Z6161: MUXCY_L port map (
    DI => R1IN_1FF(19),
    CI => R1IN_ADD_2_CRY_1,
    S => R1IN_ADD_2_AXB_2,
    LO => R1IN_ADD_2_CRY_2);
R1IN_ADD_2_S_1: XORCY port map (
    LI => R1IN_ADD_2_AXB_1,
    CI => R1IN_ADD_2_CRY_0,
    O => PRODUCT(18));
R1IN_ADD_2_CRY_1_Z6163: MUXCY_L port map (
    DI => R1IN_1FF(18),
    CI => R1IN_ADD_2_CRY_0,
    S => R1IN_ADD_2_AXB_1,
    LO => R1IN_ADD_2_CRY_1);
R1IN_ADD_2_CRY_0_Z6164: MUXCY_L port map (
    DI => R1IN_ADD_2,
    CI => NN_1,
    S => NN_3,
    LO => R1IN_ADD_2_CRY_0);
R1IN_4_4_ADD_2_S_36: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_36,
    CI => R1IN_4_4_ADD_2_CRY_35,
    O => R1IN_4_4(53));
R1IN_4_4_ADD_2_S_35: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_35,
    CI => R1IN_4_4_ADD_2_CRY_34,
    O => R1IN_4_4(52));
R1IN_4_4_ADD_2_CRY_35_Z6167: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_4_ADD_2_CRY_34,
    S => R1IN_4_4_ADD_2_AXB_35,
    LO => R1IN_4_4_ADD_2_CRY_35);
R1IN_4_4_ADD_2_S_34: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_34,
    CI => R1IN_4_4_ADD_2_CRY_33,
    O => R1IN_4_4(51));
R1IN_4_4_ADD_2_CRY_34_Z6169: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_4_ADD_2_CRY_33,
    S => R1IN_4_4_ADD_2_AXB_34,
    LO => R1IN_4_4_ADD_2_CRY_34);
R1IN_4_4_ADD_2_S_33: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_33,
    CI => R1IN_4_4_ADD_2_CRY_32,
    O => R1IN_4_4(50));
R1IN_4_4_ADD_2_CRY_33_Z6171: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_4_ADD_2_CRY_32,
    S => R1IN_4_4_ADD_2_AXB_33,
    LO => R1IN_4_4_ADD_2_CRY_33);
R1IN_4_4_ADD_2_S_32: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_32,
    CI => R1IN_4_4_ADD_2_CRY_31,
    O => R1IN_4_4(49));
R1IN_4_4_ADD_2_CRY_32_Z6173: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_4_ADD_2_CRY_31,
    S => R1IN_4_4_ADD_2_AXB_32,
    LO => R1IN_4_4_ADD_2_CRY_32);
R1IN_4_4_ADD_2_S_31: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_31,
    CI => R1IN_4_4_ADD_2_CRY_30,
    O => R1IN_4_4(48));
R1IN_4_4_ADD_2_CRY_31_Z6175: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_4_ADD_2_CRY_30,
    S => R1IN_4_4_ADD_2_AXB_31,
    LO => R1IN_4_4_ADD_2_CRY_31);
R1IN_4_4_ADD_2_S_30: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_30,
    CI => R1IN_4_4_ADD_2_CRY_29,
    O => R1IN_4_4(47));
R1IN_4_4_ADD_2_CRY_30_Z6177: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_4_ADD_2_CRY_29,
    S => R1IN_4_4_ADD_2_AXB_30,
    LO => R1IN_4_4_ADD_2_CRY_30);
R1IN_4_4_ADD_2_S_29: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_29,
    CI => R1IN_4_4_ADD_2_CRY_28,
    O => R1IN_4_4(46));
R1IN_4_4_ADD_2_CRY_29_Z6179: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_4_ADD_2_CRY_28,
    S => R1IN_4_4_ADD_2_AXB_29,
    LO => R1IN_4_4_ADD_2_CRY_29);
R1IN_4_4_ADD_2_S_28: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_28,
    CI => R1IN_4_4_ADD_2_CRY_27,
    O => R1IN_4_4(45));
R1IN_4_4_ADD_2_CRY_28_Z6181: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_4_ADD_2_CRY_27,
    S => R1IN_4_4_ADD_2_AXB_28,
    LO => R1IN_4_4_ADD_2_CRY_28);
R1IN_4_4_ADD_2_S_27: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_27,
    CI => R1IN_4_4_ADD_2_CRY_26,
    O => R1IN_4_4(44));
R1IN_4_4_ADD_2_CRY_27_Z6183: MUXCY_L port map (
    DI => R1IN_4_4_4F_RETO(10),
    CI => R1IN_4_4_ADD_2_CRY_26,
    S => R1IN_4_4_ADD_2_AXB_27,
    LO => R1IN_4_4_ADD_2_CRY_27);
R1IN_4_4_ADD_2_S_26: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_26,
    CI => R1IN_4_4_ADD_2_CRY_25,
    O => R1IN_4_4(43));
R1IN_4_4_ADD_2_CRY_26_Z6185: MUXCY_L port map (
    DI => R1IN_4_4_4F_RETO(9),
    CI => R1IN_4_4_ADD_2_CRY_25,
    S => R1IN_4_4_ADD_2_AXB_26,
    LO => R1IN_4_4_ADD_2_CRY_26);
R1IN_4_4_ADD_2_S_25: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_25,
    CI => R1IN_4_4_ADD_2_CRY_24,
    O => R1IN_4_4(42));
R1IN_4_4_ADD_2_CRY_25_Z6187: MUXCY_L port map (
    DI => R1IN_4_4_4F_RETO(8),
    CI => R1IN_4_4_ADD_2_CRY_24,
    S => R1IN_4_4_ADD_2_AXB_25,
    LO => R1IN_4_4_ADD_2_CRY_25);
R1IN_4_4_ADD_2_S_24: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_24,
    CI => R1IN_4_4_ADD_2_CRY_23,
    O => R1IN_4_4(41));
R1IN_4_4_ADD_2_CRY_24_Z6189: MUXCY_L port map (
    DI => R1IN_4_4_4F_RETO(7),
    CI => R1IN_4_4_ADD_2_CRY_23,
    S => R1IN_4_4_ADD_2_AXB_24,
    LO => R1IN_4_4_ADD_2_CRY_24);
R1IN_4_4_ADD_2_S_23: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_23,
    CI => R1IN_4_4_ADD_2_CRY_22,
    O => R1IN_4_4(40));
R1IN_4_4_ADD_2_CRY_23_Z6191: MUXCY_L port map (
    DI => R1IN_4_4_4F_RETO(6),
    CI => R1IN_4_4_ADD_2_CRY_22,
    S => R1IN_4_4_ADD_2_AXB_23,
    LO => R1IN_4_4_ADD_2_CRY_23);
R1IN_4_4_ADD_2_S_22: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_22,
    CI => R1IN_4_4_ADD_2_CRY_21,
    O => R1IN_4_4(39));
R1IN_4_4_ADD_2_CRY_22_Z6193: MUXCY_L port map (
    DI => R1IN_4_4_4F_RETO(5),
    CI => R1IN_4_4_ADD_2_CRY_21,
    S => R1IN_4_4_ADD_2_AXB_22,
    LO => R1IN_4_4_ADD_2_CRY_22);
R1IN_4_4_ADD_2_S_21: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_21,
    CI => R1IN_4_4_ADD_2_CRY_20,
    O => R1IN_4_4(38));
R1IN_4_4_ADD_2_CRY_21_Z6195: MUXCY_L port map (
    DI => R1IN_4_4_4F_RETO(4),
    CI => R1IN_4_4_ADD_2_CRY_20,
    S => R1IN_4_4_ADD_2_AXB_21,
    LO => R1IN_4_4_ADD_2_CRY_21);
R1IN_4_4_ADD_2_S_20: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_20,
    CI => R1IN_4_4_ADD_2_CRY_19,
    O => R1IN_4_4(37));
R1IN_4_4_ADD_2_CRY_20_Z6197: MUXCY_L port map (
    DI => R1IN_4_4_4F_RETO(3),
    CI => R1IN_4_4_ADD_2_CRY_19,
    S => R1IN_4_4_ADD_2_AXB_20,
    LO => R1IN_4_4_ADD_2_CRY_20);
R1IN_4_4_ADD_2_S_19: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_19,
    CI => R1IN_4_4_ADD_2_CRY_18,
    O => R1IN_4_4(36));
R1IN_4_4_ADD_2_CRY_19_Z6199: MUXCY_L port map (
    DI => R1IN_4_4_4F_RETO(2),
    CI => R1IN_4_4_ADD_2_CRY_18,
    S => R1IN_4_4_ADD_2_AXB_19,
    LO => R1IN_4_4_ADD_2_CRY_19);
R1IN_4_4_ADD_2_S_18: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_18,
    CI => R1IN_4_4_ADD_2_CRY_17,
    O => R1IN_4_4(35));
R1IN_4_4_ADD_2_CRY_18_Z6201: MUXCY_L port map (
    DI => R1IN_4_4_4F_RETO(1),
    CI => R1IN_4_4_ADD_2_CRY_17,
    S => R1IN_4_4_ADD_2_AXB_18,
    LO => R1IN_4_4_ADD_2_CRY_18);
R1IN_4_4_ADD_2_S_17: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_17,
    CI => R1IN_4_4_ADD_2_CRY_16,
    O => R1IN_4_4(34));
R1IN_4_4_ADD_2_CRY_17_Z6203: MUXCY_L port map (
    DI => R1IN_4_4_4F_RETO(0),
    CI => R1IN_4_4_ADD_2_CRY_16,
    S => R1IN_4_4_ADD_2_AXB_17,
    LO => R1IN_4_4_ADD_2_CRY_17);
R1IN_4_4_ADD_2_S_16: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_16,
    CI => R1IN_4_4_ADD_2_CRY_15,
    O => R1IN_4_4(33));
R1IN_4_4_ADD_2_CRY_16_Z6205: MUXCY_L port map (
    DI => R1IN_4_4_1F_RETO(33),
    CI => R1IN_4_4_ADD_2_CRY_15,
    S => R1IN_4_4_ADD_2_AXB_16,
    LO => R1IN_4_4_ADD_2_CRY_16);
R1IN_4_4_ADD_2_S_15: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_15,
    CI => R1IN_4_4_ADD_2_CRY_14,
    O => R1IN_4_4(32));
R1IN_4_4_ADD_2_CRY_15_Z6207: MUXCY_L port map (
    DI => R1IN_4_4_1F_RETO(32),
    CI => R1IN_4_4_ADD_2_CRY_14,
    S => R1IN_4_4_ADD_2_AXB_15,
    LO => R1IN_4_4_ADD_2_CRY_15);
R1IN_4_4_ADD_2_S_14: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_14,
    CI => R1IN_4_4_ADD_2_CRY_13,
    O => R1IN_4_4(31));
R1IN_4_4_ADD_2_CRY_14_Z6209: MUXCY_L port map (
    DI => R1IN_4_4_1F_RETO(31),
    CI => R1IN_4_4_ADD_2_CRY_13,
    S => R1IN_4_4_ADD_2_AXB_14,
    LO => R1IN_4_4_ADD_2_CRY_14);
R1IN_4_4_ADD_2_S_13: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_13,
    CI => R1IN_4_4_ADD_2_CRY_12,
    O => R1IN_4_4(30));
R1IN_4_4_ADD_2_CRY_13_Z6211: MUXCY_L port map (
    DI => R1IN_4_4_1F_RETO(30),
    CI => R1IN_4_4_ADD_2_CRY_12,
    S => R1IN_4_4_ADD_2_AXB_13,
    LO => R1IN_4_4_ADD_2_CRY_13);
R1IN_4_4_ADD_2_S_12: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_12,
    CI => R1IN_4_4_ADD_2_CRY_11,
    O => R1IN_4_4(29));
R1IN_4_4_ADD_2_CRY_12_Z6213: MUXCY_L port map (
    DI => R1IN_4_4_1F_RETO(29),
    CI => R1IN_4_4_ADD_2_CRY_11,
    S => R1IN_4_4_ADD_2_AXB_12,
    LO => R1IN_4_4_ADD_2_CRY_12);
R1IN_4_4_ADD_2_S_11: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_11,
    CI => R1IN_4_4_ADD_2_CRY_10,
    O => R1IN_4_4(28));
R1IN_4_4_ADD_2_CRY_11_Z6215: MUXCY_L port map (
    DI => R1IN_4_4_1F_RETO(28),
    CI => R1IN_4_4_ADD_2_CRY_10,
    S => R1IN_4_4_ADD_2_AXB_11,
    LO => R1IN_4_4_ADD_2_CRY_11);
R1IN_4_4_ADD_2_S_10: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_10,
    CI => R1IN_4_4_ADD_2_CRY_9,
    O => R1IN_4_4(27));
R1IN_4_4_ADD_2_CRY_10_Z6217: MUXCY_L port map (
    DI => R1IN_4_4_1F_RETO(27),
    CI => R1IN_4_4_ADD_2_CRY_9,
    S => R1IN_4_4_ADD_2_AXB_10,
    LO => R1IN_4_4_ADD_2_CRY_10);
R1IN_4_4_ADD_2_S_9: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_9,
    CI => R1IN_4_4_ADD_2_CRY_8,
    O => R1IN_4_4(26));
R1IN_4_4_ADD_2_CRY_9_Z6219: MUXCY_L port map (
    DI => R1IN_4_4_1F_RETO(26),
    CI => R1IN_4_4_ADD_2_CRY_8,
    S => R1IN_4_4_ADD_2_AXB_9,
    LO => R1IN_4_4_ADD_2_CRY_9);
R1IN_4_4_ADD_2_S_8: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_8,
    CI => R1IN_4_4_ADD_2_CRY_7,
    O => R1IN_4_4(25));
R1IN_4_4_ADD_2_CRY_8_Z6221: MUXCY_L port map (
    DI => R1IN_4_4_1F_RETO(25),
    CI => R1IN_4_4_ADD_2_CRY_7,
    S => R1IN_4_4_ADD_2_AXB_8,
    LO => R1IN_4_4_ADD_2_CRY_8);
R1IN_4_4_ADD_2_S_7: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_7,
    CI => R1IN_4_4_ADD_2_CRY_6,
    O => R1IN_4_4(24));
R1IN_4_4_ADD_2_CRY_7_Z6223: MUXCY_L port map (
    DI => R1IN_4_4_1F_RETO(24),
    CI => R1IN_4_4_ADD_2_CRY_6,
    S => R1IN_4_4_ADD_2_AXB_7,
    LO => R1IN_4_4_ADD_2_CRY_7);
R1IN_4_4_ADD_2_S_6: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_6,
    CI => R1IN_4_4_ADD_2_CRY_5,
    O => R1IN_4_4(23));
R1IN_4_4_ADD_2_CRY_6_Z6225: MUXCY_L port map (
    DI => R1IN_4_4_1F_RETO(23),
    CI => R1IN_4_4_ADD_2_CRY_5,
    S => R1IN_4_4_ADD_2_AXB_6,
    LO => R1IN_4_4_ADD_2_CRY_6);
R1IN_4_4_ADD_2_S_5: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_5,
    CI => R1IN_4_4_ADD_2_CRY_4,
    O => R1IN_4_4(22));
R1IN_4_4_ADD_2_CRY_5_Z6227: MUXCY_L port map (
    DI => R1IN_4_4_1F_RETO(22),
    CI => R1IN_4_4_ADD_2_CRY_4,
    S => R1IN_4_4_ADD_2_AXB_5,
    LO => R1IN_4_4_ADD_2_CRY_5);
R1IN_4_4_ADD_2_S_4: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_4,
    CI => R1IN_4_4_ADD_2_CRY_3,
    O => R1IN_4_4(21));
R1IN_4_4_ADD_2_CRY_4_Z6229: MUXCY_L port map (
    DI => R1IN_4_4_1F_RETO(21),
    CI => R1IN_4_4_ADD_2_CRY_3,
    S => R1IN_4_4_ADD_2_AXB_4,
    LO => R1IN_4_4_ADD_2_CRY_4);
R1IN_4_4_ADD_2_S_3: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_3,
    CI => R1IN_4_4_ADD_2_CRY_2,
    O => R1IN_4_4(20));
R1IN_4_4_ADD_2_CRY_3_Z6231: MUXCY_L port map (
    DI => R1IN_4_4_1F_RETO(20),
    CI => R1IN_4_4_ADD_2_CRY_2,
    S => R1IN_4_4_ADD_2_AXB_3,
    LO => R1IN_4_4_ADD_2_CRY_3);
R1IN_4_4_ADD_2_S_2: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_2,
    CI => R1IN_4_4_ADD_2_CRY_1,
    O => R1IN_4_4(19));
R1IN_4_4_ADD_2_CRY_2_Z6233: MUXCY_L port map (
    DI => R1IN_4_4_1F_RETO(19),
    CI => R1IN_4_4_ADD_2_CRY_1,
    S => R1IN_4_4_ADD_2_AXB_2,
    LO => R1IN_4_4_ADD_2_CRY_2);
R1IN_4_4_ADD_2_S_1: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_1,
    CI => R1IN_4_4_ADD_2_CRY_0,
    O => R1IN_4_4(18));
R1IN_4_4_ADD_2_CRY_1_Z6235: MUXCY_L port map (
    DI => R1IN_4_4_1F_RETO(18),
    CI => R1IN_4_4_ADD_2_CRY_0,
    S => R1IN_4_4_ADD_2_AXB_1,
    LO => R1IN_4_4_ADD_2_CRY_1);
R1IN_4_4_ADD_2_CRY_0_Z6236: MUXCY_L port map (
    DI => R1IN_4_4_ADD_2_RETO_0,
    CI => NN_1,
    S => R1IN_4_4(17),
    LO => R1IN_4_4_ADD_2_CRY_0);
R1IN_3_ADD_1_S_43: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_43,
    CI => R1IN_3_ADD_1_CRY_42,
    O => R1IN_3(60));
R1IN_3_ADD_1_S_42: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_42,
    CI => R1IN_3_ADD_1_CRY_41,
    O => R1IN_3(59));
R1IN_3_ADD_1_CRY_42_Z6239: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_41,
    S => R1IN_3_ADD_1_AXB_42,
    LO => R1IN_3_ADD_1_CRY_42);
R1IN_3_ADD_1_S_41: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_41,
    CI => R1IN_3_ADD_1_CRY_40,
    O => R1IN_3(58));
R1IN_3_ADD_1_CRY_41_Z6241: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_40,
    S => R1IN_3_ADD_1_AXB_41,
    LO => R1IN_3_ADD_1_CRY_41);
R1IN_3_ADD_1_S_40: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_40,
    CI => R1IN_3_ADD_1_CRY_39,
    O => R1IN_3(57));
R1IN_3_ADD_1_CRY_40_Z6243: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_39,
    S => R1IN_3_ADD_1_AXB_40,
    LO => R1IN_3_ADD_1_CRY_40);
R1IN_3_ADD_1_S_39: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_39,
    CI => R1IN_3_ADD_1_CRY_38,
    O => R1IN_3(56));
R1IN_3_ADD_1_CRY_39_Z6245: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_38,
    S => R1IN_3_ADD_1_AXB_39,
    LO => R1IN_3_ADD_1_CRY_39);
R1IN_3_ADD_1_S_38: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_38,
    CI => R1IN_3_ADD_1_CRY_37,
    O => R1IN_3(55));
R1IN_3_ADD_1_CRY_38_Z6247: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_37,
    S => R1IN_3_ADD_1_AXB_38,
    LO => R1IN_3_ADD_1_CRY_38);
R1IN_3_ADD_1_S_37: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_37,
    CI => R1IN_3_ADD_1_CRY_36,
    O => R1IN_3(54));
R1IN_3_ADD_1_CRY_37_Z6249: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_36,
    S => R1IN_3_ADD_1_AXB_37,
    LO => R1IN_3_ADD_1_CRY_37);
R1IN_3_ADD_1_S_36: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_36,
    CI => R1IN_3_ADD_1_CRY_35,
    O => R1IN_3(53));
R1IN_3_ADD_1_CRY_36_Z6251: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_35,
    S => R1IN_3_ADD_1_AXB_36,
    LO => R1IN_3_ADD_1_CRY_36);
R1IN_3_ADD_1_S_35: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_35,
    CI => R1IN_3_ADD_1_CRY_34,
    O => R1IN_3(52));
R1IN_3_ADD_1_CRY_35_Z6253: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_34,
    S => R1IN_3_ADD_1_AXB_35,
    LO => R1IN_3_ADD_1_CRY_35);
R1IN_3_ADD_1_S_34: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_34,
    CI => R1IN_3_ADD_1_CRY_33,
    O => R1IN_3(51));
R1IN_3_ADD_1_CRY_34_Z6255: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_33,
    S => R1IN_3_ADD_1_AXB_34,
    LO => R1IN_3_ADD_1_CRY_34);
R1IN_3_ADD_1_S_33: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_33,
    CI => R1IN_3_ADD_1_CRY_32,
    O => R1IN_3(50));
R1IN_3_ADD_1_CRY_33_Z6257: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_32,
    S => R1IN_3_ADD_1_AXB_33,
    LO => R1IN_3_ADD_1_CRY_33);
R1IN_3_ADD_1_S_32: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_32,
    CI => R1IN_3_ADD_1_CRY_31,
    O => R1IN_3(49));
R1IN_3_ADD_1_CRY_32_Z6259: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_31,
    S => R1IN_3_ADD_1_AXB_32,
    LO => R1IN_3_ADD_1_CRY_32);
R1IN_3_ADD_1_S_31: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_31,
    CI => R1IN_3_ADD_1_CRY_30,
    O => R1IN_3(48));
R1IN_3_ADD_1_CRY_31_Z6261: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_30,
    S => R1IN_3_ADD_1_AXB_31,
    LO => R1IN_3_ADD_1_CRY_31);
R1IN_3_ADD_1_S_30: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_30,
    CI => R1IN_3_ADD_1_CRY_29,
    O => R1IN_3(47));
R1IN_3_ADD_1_CRY_30_Z6263: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_29,
    S => R1IN_3_ADD_1_AXB_30,
    LO => R1IN_3_ADD_1_CRY_30);
R1IN_3_ADD_1_S_29: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_29,
    CI => R1IN_3_ADD_1_CRY_28,
    O => R1IN_3(46));
R1IN_3_ADD_1_CRY_29_Z6265: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_28,
    S => R1IN_3_ADD_1_AXB_29,
    LO => R1IN_3_ADD_1_CRY_29);
R1IN_3_ADD_1_S_28: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_28,
    CI => R1IN_3_ADD_1_CRY_27,
    O => R1IN_3(45));
R1IN_3_ADD_1_CRY_28_Z6267: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_27,
    S => R1IN_3_ADD_1_AXB_28,
    LO => R1IN_3_ADD_1_CRY_28);
R1IN_3_ADD_1_S_27: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_27,
    CI => R1IN_3_ADD_1_CRY_26,
    O => R1IN_3(44));
R1IN_3_ADD_1_CRY_27_Z6269: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_26,
    S => R1IN_3_ADD_1_AXB_27,
    LO => R1IN_3_ADD_1_CRY_27);
R1IN_3_ADD_1_S_26: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_26,
    CI => R1IN_3_ADD_1_CRY_25,
    O => R1IN_3(43));
R1IN_3_ADD_1_CRY_26_Z6271: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_25,
    S => R1IN_3_ADD_1_AXB_26,
    LO => R1IN_3_ADD_1_CRY_26);
R1IN_3_ADD_1_S_25: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_25,
    CI => R1IN_3_ADD_1_CRY_24,
    O => R1IN_3(42));
R1IN_3_ADD_1_CRY_25_Z6273: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_24,
    S => R1IN_3_ADD_1_AXB_25,
    LO => R1IN_3_ADD_1_CRY_25);
R1IN_3_ADD_1_S_24: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_24,
    CI => R1IN_3_ADD_1_CRY_23,
    O => R1IN_3(41));
R1IN_3_ADD_1_CRY_24_Z6275: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_23,
    S => R1IN_3_ADD_1_AXB_24,
    LO => R1IN_3_ADD_1_CRY_24);
R1IN_3_ADD_1_S_23: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_23,
    CI => R1IN_3_ADD_1_CRY_22,
    O => R1IN_3(40));
R1IN_3_ADD_1_CRY_23_Z6277: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_22,
    S => R1IN_3_ADD_1_AXB_23,
    LO => R1IN_3_ADD_1_CRY_23);
R1IN_3_ADD_1_S_22: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_22,
    CI => R1IN_3_ADD_1_CRY_21,
    O => R1IN_3(39));
R1IN_3_ADD_1_CRY_22_Z6279: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_21,
    S => R1IN_3_ADD_1_AXB_22,
    LO => R1IN_3_ADD_1_CRY_22);
R1IN_3_ADD_1_S_21: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_21,
    CI => R1IN_3_ADD_1_CRY_20,
    O => R1IN_3(38));
R1IN_3_ADD_1_CRY_21_Z6281: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_20,
    S => R1IN_3_ADD_1_AXB_21,
    LO => R1IN_3_ADD_1_CRY_21);
R1IN_3_ADD_1_S_20: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_20,
    CI => R1IN_3_ADD_1_CRY_19,
    O => R1IN_3(37));
R1IN_3_ADD_1_CRY_20_Z6283: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_19,
    S => R1IN_3_ADD_1_AXB_20,
    LO => R1IN_3_ADD_1_CRY_20);
R1IN_3_ADD_1_S_19: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_19,
    CI => R1IN_3_ADD_1_CRY_18,
    O => R1IN_3(36));
R1IN_3_ADD_1_CRY_19_Z6285: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_18,
    S => R1IN_3_ADD_1_AXB_19,
    LO => R1IN_3_ADD_1_CRY_19);
R1IN_3_ADD_1_S_18: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_18,
    CI => R1IN_3_ADD_1_CRY_17,
    O => R1IN_3(35));
R1IN_3_ADD_1_CRY_18_Z6287: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_17,
    S => R1IN_3_ADD_1_AXB_18,
    LO => R1IN_3_ADD_1_CRY_18);
R1IN_3_ADD_1_S_17: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_17,
    CI => R1IN_3_ADD_1_CRY_16,
    O => R1IN_3(34));
R1IN_3_ADD_1_CRY_17_Z6289: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_16,
    S => R1IN_3_ADD_1_AXB_17,
    LO => R1IN_3_ADD_1_CRY_17);
R1IN_3_ADD_1_S_16: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_16,
    CI => R1IN_3_ADD_1_CRY_15,
    O => R1IN_3(33));
R1IN_3_ADD_1_CRY_16_Z6291: MUXCY_L port map (
    DI => R1IN_3_2F_RETO(16),
    CI => R1IN_3_ADD_1_CRY_15,
    S => R1IN_3_ADD_1_AXB_16,
    LO => R1IN_3_ADD_1_CRY_16);
R1IN_3_ADD_1_S_15: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_15,
    CI => R1IN_3_ADD_1_CRY_14,
    O => R1IN_3(32));
R1IN_3_ADD_1_CRY_15_Z6293: MUXCY_L port map (
    DI => R1IN_3_2F_RETO(15),
    CI => R1IN_3_ADD_1_CRY_14,
    S => R1IN_3_ADD_1_AXB_15,
    LO => R1IN_3_ADD_1_CRY_15);
R1IN_3_ADD_1_S_14: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_14,
    CI => R1IN_3_ADD_1_CRY_13,
    O => R1IN_3(31));
R1IN_3_ADD_1_CRY_14_Z6295: MUXCY_L port map (
    DI => R1IN_3_2F_RETO(14),
    CI => R1IN_3_ADD_1_CRY_13,
    S => R1IN_3_ADD_1_AXB_14,
    LO => R1IN_3_ADD_1_CRY_14);
R1IN_3_ADD_1_S_13: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_13,
    CI => R1IN_3_ADD_1_CRY_12,
    O => R1IN_3(30));
R1IN_3_ADD_1_CRY_13_Z6297: MUXCY_L port map (
    DI => R1IN_3_2F_RETO(13),
    CI => R1IN_3_ADD_1_CRY_12,
    S => R1IN_3_ADD_1_AXB_13,
    LO => R1IN_3_ADD_1_CRY_13);
R1IN_3_ADD_1_S_12: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_12,
    CI => R1IN_3_ADD_1_CRY_11,
    O => R1IN_3(29));
R1IN_3_ADD_1_CRY_12_Z6299: MUXCY_L port map (
    DI => R1IN_3_2F_RETO(12),
    CI => R1IN_3_ADD_1_CRY_11,
    S => R1IN_3_ADD_1_AXB_12,
    LO => R1IN_3_ADD_1_CRY_12);
R1IN_3_ADD_1_S_11: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_11,
    CI => R1IN_3_ADD_1_CRY_10,
    O => R1IN_3(28));
R1IN_3_ADD_1_CRY_11_Z6301: MUXCY_L port map (
    DI => R1IN_3_2F_RETO(11),
    CI => R1IN_3_ADD_1_CRY_10,
    S => R1IN_3_ADD_1_AXB_11,
    LO => R1IN_3_ADD_1_CRY_11);
R1IN_3_ADD_1_S_10: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_10,
    CI => R1IN_3_ADD_1_CRY_9,
    O => R1IN_3(27));
R1IN_3_ADD_1_CRY_10_Z6303: MUXCY_L port map (
    DI => R1IN_3_2F_RETO(10),
    CI => R1IN_3_ADD_1_CRY_9,
    S => R1IN_3_ADD_1_AXB_10,
    LO => R1IN_3_ADD_1_CRY_10);
R1IN_3_ADD_1_S_9: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_9,
    CI => R1IN_3_ADD_1_CRY_8,
    O => R1IN_3(26));
R1IN_3_ADD_1_CRY_9_Z6305: MUXCY_L port map (
    DI => R1IN_3_2F_RETO(9),
    CI => R1IN_3_ADD_1_CRY_8,
    S => R1IN_3_ADD_1_AXB_9,
    LO => R1IN_3_ADD_1_CRY_9);
R1IN_3_ADD_1_S_8: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_8,
    CI => R1IN_3_ADD_1_CRY_7,
    O => R1IN_3(25));
R1IN_3_ADD_1_CRY_8_Z6307: MUXCY_L port map (
    DI => R1IN_3_2F_RETO(8),
    CI => R1IN_3_ADD_1_CRY_7,
    S => R1IN_3_ADD_1_AXB_8,
    LO => R1IN_3_ADD_1_CRY_8);
R1IN_3_ADD_1_S_7: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_7,
    CI => R1IN_3_ADD_1_CRY_6,
    O => R1IN_3(24));
R1IN_3_ADD_1_CRY_7_Z6309: MUXCY_L port map (
    DI => R1IN_3_2F_RETO(7),
    CI => R1IN_3_ADD_1_CRY_6,
    S => R1IN_3_ADD_1_AXB_7,
    LO => R1IN_3_ADD_1_CRY_7);
R1IN_3_ADD_1_S_6: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_6,
    CI => R1IN_3_ADD_1_CRY_5,
    O => R1IN_3(23));
R1IN_3_ADD_1_CRY_6_Z6311: MUXCY_L port map (
    DI => R1IN_3_2F_RETO(6),
    CI => R1IN_3_ADD_1_CRY_5,
    S => R1IN_3_ADD_1_AXB_6,
    LO => R1IN_3_ADD_1_CRY_6);
R1IN_3_ADD_1_S_5: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_5,
    CI => R1IN_3_ADD_1_CRY_4,
    O => R1IN_3(22));
R1IN_3_ADD_1_CRY_5_Z6313: MUXCY_L port map (
    DI => R1IN_3_2F_RETO(5),
    CI => R1IN_3_ADD_1_CRY_4,
    S => R1IN_3_ADD_1_AXB_5,
    LO => R1IN_3_ADD_1_CRY_5);
R1IN_3_ADD_1_S_4: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_4,
    CI => R1IN_3_ADD_1_CRY_3,
    O => R1IN_3(21));
R1IN_3_ADD_1_CRY_4_Z6315: MUXCY_L port map (
    DI => R1IN_3_2F_RETO(4),
    CI => R1IN_3_ADD_1_CRY_3,
    S => R1IN_3_ADD_1_AXB_4,
    LO => R1IN_3_ADD_1_CRY_4);
R1IN_3_ADD_1_S_3: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_3,
    CI => R1IN_3_ADD_1_CRY_2,
    O => R1IN_3(20));
R1IN_3_ADD_1_CRY_3_Z6317: MUXCY_L port map (
    DI => R1IN_3_2F_RETO(3),
    CI => R1IN_3_ADD_1_CRY_2,
    S => R1IN_3_ADD_1_AXB_3,
    LO => R1IN_3_ADD_1_CRY_3);
R1IN_3_ADD_1_S_2: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_2,
    CI => R1IN_3_ADD_1_CRY_1,
    O => R1IN_3(19));
R1IN_3_ADD_1_CRY_2_Z6319: MUXCY_L port map (
    DI => R1IN_3_2F_RETO(2),
    CI => R1IN_3_ADD_1_CRY_1,
    S => R1IN_3_ADD_1_AXB_2,
    LO => R1IN_3_ADD_1_CRY_2);
R1IN_3_ADD_1_S_1: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_1,
    CI => R1IN_3_ADD_1_CRY_0,
    O => R1IN_3(18));
R1IN_3_ADD_1_CRY_1_Z6321: MUXCY_L port map (
    DI => R1IN_3_2F_RETO(1),
    CI => R1IN_3_ADD_1_CRY_0,
    S => R1IN_3_ADD_1_AXB_1,
    LO => R1IN_3_ADD_1_CRY_1);
R1IN_3_ADD_1_CRY_0_Z6322: MUXCY_L port map (
    DI => R1IN_3_ADD_1_RETO_0,
    CI => NN_1,
    S => R1IN_3(17),
    LO => R1IN_3_ADD_1_CRY_0);
R1IN_ADD_1_1_0_S_28: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_28,
    CI => R1IN_ADD_1_1_0_CRY_27,
    O => N_1592);
R1IN_ADD_1_1_0_CRY_28_Z6324: MUXCY port map (
    DI => R1IN_3(60),
    CI => R1IN_ADD_1_1_0_CRY_27,
    S => R1IN_ADD_1_1_0_AXB_28,
    O => R1IN_ADD_1_1_0_CRY_28);
R1IN_ADD_1_1_0_S_27: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_27,
    CI => R1IN_ADD_1_1_0_CRY_26,
    O => N_1591);
R1IN_ADD_1_1_0_CRY_27_Z6326: MUXCY_L port map (
    DI => R1IN_3(59),
    CI => R1IN_ADD_1_1_0_CRY_26,
    S => R1IN_ADD_1_1_0_AXB_27,
    LO => R1IN_ADD_1_1_0_CRY_27);
R1IN_ADD_1_1_0_S_26: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_26,
    CI => R1IN_ADD_1_1_0_CRY_25,
    O => N_1590);
R1IN_ADD_1_1_0_CRY_26_Z6328: MUXCY_L port map (
    DI => R1IN_3(58),
    CI => R1IN_ADD_1_1_0_CRY_25,
    S => R1IN_ADD_1_1_0_AXB_26,
    LO => R1IN_ADD_1_1_0_CRY_26);
R1IN_ADD_1_1_0_S_25: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_25,
    CI => R1IN_ADD_1_1_0_CRY_24,
    O => N_1589);
R1IN_ADD_1_1_0_CRY_25_Z6330: MUXCY_L port map (
    DI => R1IN_3(57),
    CI => R1IN_ADD_1_1_0_CRY_24,
    S => R1IN_ADD_1_1_0_AXB_25,
    LO => R1IN_ADD_1_1_0_CRY_25);
R1IN_ADD_1_1_0_S_24: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_24,
    CI => R1IN_ADD_1_1_0_CRY_23,
    O => N_1588);
R1IN_ADD_1_1_0_CRY_24_Z6332: MUXCY_L port map (
    DI => R1IN_3(56),
    CI => R1IN_ADD_1_1_0_CRY_23,
    S => R1IN_ADD_1_1_0_AXB_24,
    LO => R1IN_ADD_1_1_0_CRY_24);
R1IN_ADD_1_1_0_S_23: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_23,
    CI => R1IN_ADD_1_1_0_CRY_22,
    O => N_1587);
R1IN_ADD_1_1_0_CRY_23_Z6334: MUXCY_L port map (
    DI => R1IN_3(55),
    CI => R1IN_ADD_1_1_0_CRY_22,
    S => R1IN_ADD_1_1_0_AXB_23,
    LO => R1IN_ADD_1_1_0_CRY_23);
R1IN_ADD_1_1_0_S_22: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_22,
    CI => R1IN_ADD_1_1_0_CRY_21,
    O => N_1586);
R1IN_ADD_1_1_0_CRY_22_Z6336: MUXCY_L port map (
    DI => R1IN_3(54),
    CI => R1IN_ADD_1_1_0_CRY_21,
    S => R1IN_ADD_1_1_0_AXB_22,
    LO => R1IN_ADD_1_1_0_CRY_22);
R1IN_ADD_1_1_0_S_21: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_21,
    CI => R1IN_ADD_1_1_0_CRY_20,
    O => N_1585);
R1IN_ADD_1_1_0_CRY_21_Z6338: MUXCY_L port map (
    DI => R1IN_3(53),
    CI => R1IN_ADD_1_1_0_CRY_20,
    S => R1IN_ADD_1_1_0_AXB_21,
    LO => R1IN_ADD_1_1_0_CRY_21);
R1IN_ADD_1_1_0_S_20: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_20,
    CI => R1IN_ADD_1_1_0_CRY_19,
    O => N_1584);
R1IN_ADD_1_1_0_CRY_20_Z6340: MUXCY_L port map (
    DI => R1IN_3(52),
    CI => R1IN_ADD_1_1_0_CRY_19,
    S => R1IN_ADD_1_1_0_AXB_20,
    LO => R1IN_ADD_1_1_0_CRY_20);
R1IN_ADD_1_1_0_S_19: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_19,
    CI => R1IN_ADD_1_1_0_CRY_18,
    O => N_1583);
R1IN_ADD_1_1_0_CRY_19_Z6342: MUXCY_L port map (
    DI => R1IN_3(51),
    CI => R1IN_ADD_1_1_0_CRY_18,
    S => R1IN_ADD_1_1_0_AXB_19,
    LO => R1IN_ADD_1_1_0_CRY_19);
R1IN_ADD_1_1_0_S_18: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_18,
    CI => R1IN_ADD_1_1_0_CRY_17,
    O => N_1582);
R1IN_ADD_1_1_0_CRY_18_Z6344: MUXCY_L port map (
    DI => R1IN_3(50),
    CI => R1IN_ADD_1_1_0_CRY_17,
    S => R1IN_ADD_1_1_0_AXB_18,
    LO => R1IN_ADD_1_1_0_CRY_18);
R1IN_ADD_1_1_0_S_17: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_17,
    CI => R1IN_ADD_1_1_0_CRY_16,
    O => N_1581);
R1IN_ADD_1_1_0_CRY_17_Z6346: MUXCY_L port map (
    DI => R1IN_3(49),
    CI => R1IN_ADD_1_1_0_CRY_16,
    S => R1IN_ADD_1_1_0_AXB_17,
    LO => R1IN_ADD_1_1_0_CRY_17);
R1IN_ADD_1_1_0_S_16: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_16,
    CI => R1IN_ADD_1_1_0_CRY_15,
    O => N_1580);
R1IN_ADD_1_1_0_CRY_16_Z6348: MUXCY_L port map (
    DI => R1IN_3(48),
    CI => R1IN_ADD_1_1_0_CRY_15,
    S => R1IN_ADD_1_1_0_AXB_16,
    LO => R1IN_ADD_1_1_0_CRY_16);
R1IN_ADD_1_1_0_S_15: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_15,
    CI => R1IN_ADD_1_1_0_CRY_14,
    O => N_1579);
R1IN_ADD_1_1_0_CRY_15_Z6350: MUXCY_L port map (
    DI => R1IN_3(47),
    CI => R1IN_ADD_1_1_0_CRY_14,
    S => R1IN_ADD_1_1_0_AXB_15,
    LO => R1IN_ADD_1_1_0_CRY_15);
R1IN_ADD_1_1_0_S_14: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_14,
    CI => R1IN_ADD_1_1_0_CRY_13,
    O => N_1578);
R1IN_ADD_1_1_0_CRY_14_Z6352: MUXCY_L port map (
    DI => R1IN_3(46),
    CI => R1IN_ADD_1_1_0_CRY_13,
    S => R1IN_ADD_1_1_0_AXB_14,
    LO => R1IN_ADD_1_1_0_CRY_14);
R1IN_ADD_1_1_0_S_13: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_13,
    CI => R1IN_ADD_1_1_0_CRY_12,
    O => N_1577);
R1IN_ADD_1_1_0_CRY_13_Z6354: MUXCY_L port map (
    DI => R1IN_3(45),
    CI => R1IN_ADD_1_1_0_CRY_12,
    S => R1IN_ADD_1_1_0_AXB_13,
    LO => R1IN_ADD_1_1_0_CRY_13);
R1IN_ADD_1_1_0_S_12: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_12,
    CI => R1IN_ADD_1_1_0_CRY_11,
    O => N_1576);
R1IN_ADD_1_1_0_CRY_12_Z6356: MUXCY_L port map (
    DI => R1IN_3(44),
    CI => R1IN_ADD_1_1_0_CRY_11,
    S => R1IN_ADD_1_1_0_AXB_12,
    LO => R1IN_ADD_1_1_0_CRY_12);
R1IN_ADD_1_1_0_S_11: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_11,
    CI => R1IN_ADD_1_1_0_CRY_10,
    O => N_1575);
R1IN_ADD_1_1_0_CRY_11_Z6358: MUXCY_L port map (
    DI => R1IN_3(43),
    CI => R1IN_ADD_1_1_0_CRY_10,
    S => R1IN_ADD_1_1_0_AXB_11,
    LO => R1IN_ADD_1_1_0_CRY_11);
R1IN_ADD_1_1_0_S_10: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_10,
    CI => R1IN_ADD_1_1_0_CRY_9,
    O => N_1574);
R1IN_ADD_1_1_0_CRY_10_Z6360: MUXCY_L port map (
    DI => R1IN_3(42),
    CI => R1IN_ADD_1_1_0_CRY_9,
    S => R1IN_ADD_1_1_0_AXB_10,
    LO => R1IN_ADD_1_1_0_CRY_10);
R1IN_ADD_1_1_0_S_9: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_9,
    CI => R1IN_ADD_1_1_0_CRY_8,
    O => N_1573);
R1IN_ADD_1_1_0_CRY_9_Z6362: MUXCY_L port map (
    DI => R1IN_3(41),
    CI => R1IN_ADD_1_1_0_CRY_8,
    S => R1IN_ADD_1_1_0_AXB_9,
    LO => R1IN_ADD_1_1_0_CRY_9);
R1IN_ADD_1_1_0_S_8: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_8,
    CI => R1IN_ADD_1_1_0_CRY_7,
    O => N_1572);
R1IN_ADD_1_1_0_CRY_8_Z6364: MUXCY_L port map (
    DI => R1IN_3(40),
    CI => R1IN_ADD_1_1_0_CRY_7,
    S => R1IN_ADD_1_1_0_AXB_8,
    LO => R1IN_ADD_1_1_0_CRY_8);
R1IN_ADD_1_1_0_S_7: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_7,
    CI => R1IN_ADD_1_1_0_CRY_6,
    O => N_1571);
R1IN_ADD_1_1_0_CRY_7_Z6366: MUXCY_L port map (
    DI => R1IN_3(39),
    CI => R1IN_ADD_1_1_0_CRY_6,
    S => R1IN_ADD_1_1_0_AXB_7,
    LO => R1IN_ADD_1_1_0_CRY_7);
R1IN_ADD_1_1_0_S_6: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_6,
    CI => R1IN_ADD_1_1_0_CRY_5,
    O => N_1570);
R1IN_ADD_1_1_0_CRY_6_Z6368: MUXCY_L port map (
    DI => R1IN_3(38),
    CI => R1IN_ADD_1_1_0_CRY_5,
    S => R1IN_ADD_1_1_0_AXB_6,
    LO => R1IN_ADD_1_1_0_CRY_6);
R1IN_ADD_1_1_0_S_5: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_5,
    CI => R1IN_ADD_1_1_0_CRY_4,
    O => N_1569);
R1IN_ADD_1_1_0_CRY_5_Z6370: MUXCY_L port map (
    DI => R1IN_3(37),
    CI => R1IN_ADD_1_1_0_CRY_4,
    S => R1IN_ADD_1_1_0_AXB_5,
    LO => R1IN_ADD_1_1_0_CRY_5);
R1IN_ADD_1_1_0_S_4: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_4,
    CI => R1IN_ADD_1_1_0_CRY_3,
    O => N_1568);
R1IN_ADD_1_1_0_CRY_4_Z6372: MUXCY_L port map (
    DI => R1IN_3(36),
    CI => R1IN_ADD_1_1_0_CRY_3,
    S => R1IN_ADD_1_1_0_AXB_4,
    LO => R1IN_ADD_1_1_0_CRY_4);
R1IN_ADD_1_1_0_S_3: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_3,
    CI => R1IN_ADD_1_1_0_CRY_2,
    O => N_1567);
R1IN_ADD_1_1_0_CRY_3_Z6374: MUXCY_L port map (
    DI => R1IN_3(35),
    CI => R1IN_ADD_1_1_0_CRY_2,
    S => R1IN_ADD_1_1_0_AXB_3,
    LO => R1IN_ADD_1_1_0_CRY_3);
R1IN_ADD_1_1_0_S_2: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_2,
    CI => R1IN_ADD_1_1_0_CRY_1,
    O => N_1566);
R1IN_ADD_1_1_0_CRY_2_Z6376: MUXCY_L port map (
    DI => R1IN_3(34),
    CI => R1IN_ADD_1_1_0_CRY_1,
    S => R1IN_ADD_1_1_0_AXB_2,
    LO => R1IN_ADD_1_1_0_CRY_2);
R1IN_ADD_1_1_0_S_1: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_1,
    CI => R1IN_ADD_1_1_0_CRY_0,
    O => N_1565);
R1IN_ADD_1_1_0_CRY_1_Z6378: MUXCY_L port map (
    DI => R1IN_3(33),
    CI => R1IN_ADD_1_1_0_CRY_0,
    S => R1IN_ADD_1_1_0_AXB_1,
    LO => R1IN_ADD_1_1_0_CRY_1);
R1IN_ADD_1_1_0_CRY_0_Z6379: MUXCY_L port map (
    DI => R1IN_3(32),
    CI => NN_2,
    S => R1IN_ADD_1_1_0_AXB_0,
    LO => R1IN_ADD_1_1_0_CRY_0);
R1IN_ADD_1_1_S_28: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_28,
    CI => R1IN_ADD_1_1_CRY_27,
    O => N_1433);
R1IN_ADD_1_1_S_27: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_27,
    CI => R1IN_ADD_1_1_CRY_26,
    O => N_1431);
R1IN_ADD_1_1_CRY_27_Z6382: MUXCY_L port map (
    DI => R1IN_3(59),
    CI => R1IN_ADD_1_1_CRY_26,
    S => R1IN_ADD_1_1_AXB_27,
    LO => R1IN_ADD_1_1_CRY_27);
R1IN_ADD_1_1_S_26: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_26,
    CI => R1IN_ADD_1_1_CRY_25,
    O => N_1429);
R1IN_ADD_1_1_CRY_26_Z6384: MUXCY_L port map (
    DI => R1IN_3(58),
    CI => R1IN_ADD_1_1_CRY_25,
    S => R1IN_ADD_1_1_AXB_26,
    LO => R1IN_ADD_1_1_CRY_26);
R1IN_ADD_1_1_S_25: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_25,
    CI => R1IN_ADD_1_1_CRY_24,
    O => N_1427);
R1IN_ADD_1_1_CRY_25_Z6386: MUXCY_L port map (
    DI => R1IN_3(57),
    CI => R1IN_ADD_1_1_CRY_24,
    S => R1IN_ADD_1_1_AXB_25,
    LO => R1IN_ADD_1_1_CRY_25);
R1IN_ADD_1_1_S_24: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_24,
    CI => R1IN_ADD_1_1_CRY_23,
    O => N_1425);
R1IN_ADD_1_1_CRY_24_Z6388: MUXCY_L port map (
    DI => R1IN_3(56),
    CI => R1IN_ADD_1_1_CRY_23,
    S => R1IN_ADD_1_1_AXB_24,
    LO => R1IN_ADD_1_1_CRY_24);
R1IN_ADD_1_1_S_23: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_23,
    CI => R1IN_ADD_1_1_CRY_22,
    O => N_1423);
R1IN_ADD_1_1_CRY_23_Z6390: MUXCY_L port map (
    DI => R1IN_3(55),
    CI => R1IN_ADD_1_1_CRY_22,
    S => R1IN_ADD_1_1_AXB_23,
    LO => R1IN_ADD_1_1_CRY_23);
R1IN_ADD_1_1_S_22: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_22,
    CI => R1IN_ADD_1_1_CRY_21,
    O => N_1421);
R1IN_ADD_1_1_CRY_22_Z6392: MUXCY_L port map (
    DI => R1IN_3(54),
    CI => R1IN_ADD_1_1_CRY_21,
    S => R1IN_ADD_1_1_AXB_22,
    LO => R1IN_ADD_1_1_CRY_22);
R1IN_ADD_1_1_S_21: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_21,
    CI => R1IN_ADD_1_1_CRY_20,
    O => N_1419);
R1IN_ADD_1_1_CRY_21_Z6394: MUXCY_L port map (
    DI => R1IN_3(53),
    CI => R1IN_ADD_1_1_CRY_20,
    S => R1IN_ADD_1_1_AXB_21,
    LO => R1IN_ADD_1_1_CRY_21);
R1IN_ADD_1_1_S_20: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_20,
    CI => R1IN_ADD_1_1_CRY_19,
    O => N_1417);
R1IN_ADD_1_1_CRY_20_Z6396: MUXCY_L port map (
    DI => R1IN_3(52),
    CI => R1IN_ADD_1_1_CRY_19,
    S => R1IN_ADD_1_1_AXB_20,
    LO => R1IN_ADD_1_1_CRY_20);
R1IN_ADD_1_1_S_19: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_19,
    CI => R1IN_ADD_1_1_CRY_18,
    O => N_1415);
R1IN_ADD_1_1_CRY_19_Z6398: MUXCY_L port map (
    DI => R1IN_3(51),
    CI => R1IN_ADD_1_1_CRY_18,
    S => R1IN_ADD_1_1_AXB_19,
    LO => R1IN_ADD_1_1_CRY_19);
R1IN_ADD_1_1_S_18: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_18,
    CI => R1IN_ADD_1_1_CRY_17,
    O => N_1413);
R1IN_ADD_1_1_CRY_18_Z6400: MUXCY_L port map (
    DI => R1IN_3(50),
    CI => R1IN_ADD_1_1_CRY_17,
    S => R1IN_ADD_1_1_AXB_18,
    LO => R1IN_ADD_1_1_CRY_18);
R1IN_ADD_1_1_S_17: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_17,
    CI => R1IN_ADD_1_1_CRY_16,
    O => N_1411);
R1IN_ADD_1_1_CRY_17_Z6402: MUXCY_L port map (
    DI => R1IN_3(49),
    CI => R1IN_ADD_1_1_CRY_16,
    S => R1IN_ADD_1_1_AXB_17,
    LO => R1IN_ADD_1_1_CRY_17);
R1IN_ADD_1_1_S_16: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_16,
    CI => R1IN_ADD_1_1_CRY_15,
    O => N_1409);
R1IN_ADD_1_1_CRY_16_Z6404: MUXCY_L port map (
    DI => R1IN_3(48),
    CI => R1IN_ADD_1_1_CRY_15,
    S => R1IN_ADD_1_1_AXB_16,
    LO => R1IN_ADD_1_1_CRY_16);
R1IN_ADD_1_1_S_15: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_15,
    CI => R1IN_ADD_1_1_CRY_14,
    O => N_1407);
R1IN_ADD_1_1_CRY_15_Z6406: MUXCY_L port map (
    DI => R1IN_3(47),
    CI => R1IN_ADD_1_1_CRY_14,
    S => R1IN_ADD_1_1_AXB_15,
    LO => R1IN_ADD_1_1_CRY_15);
R1IN_ADD_1_1_S_14: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_14,
    CI => R1IN_ADD_1_1_CRY_13,
    O => N_1405);
R1IN_ADD_1_1_CRY_14_Z6408: MUXCY_L port map (
    DI => R1IN_3(46),
    CI => R1IN_ADD_1_1_CRY_13,
    S => R1IN_ADD_1_1_AXB_14,
    LO => R1IN_ADD_1_1_CRY_14);
R1IN_ADD_1_1_S_13: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_13,
    CI => R1IN_ADD_1_1_CRY_12,
    O => N_1403);
R1IN_ADD_1_1_CRY_13_Z6410: MUXCY_L port map (
    DI => R1IN_3(45),
    CI => R1IN_ADD_1_1_CRY_12,
    S => R1IN_ADD_1_1_AXB_13,
    LO => R1IN_ADD_1_1_CRY_13);
R1IN_ADD_1_1_S_12: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_12,
    CI => R1IN_ADD_1_1_CRY_11,
    O => N_1401);
R1IN_ADD_1_1_CRY_12_Z6412: MUXCY_L port map (
    DI => R1IN_3(44),
    CI => R1IN_ADD_1_1_CRY_11,
    S => R1IN_ADD_1_1_AXB_12,
    LO => R1IN_ADD_1_1_CRY_12);
R1IN_ADD_1_1_S_11: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_11,
    CI => R1IN_ADD_1_1_CRY_10,
    O => N_1399);
R1IN_ADD_1_1_CRY_11_Z6414: MUXCY_L port map (
    DI => R1IN_3(43),
    CI => R1IN_ADD_1_1_CRY_10,
    S => R1IN_ADD_1_1_AXB_11,
    LO => R1IN_ADD_1_1_CRY_11);
R1IN_ADD_1_1_S_10: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_10,
    CI => R1IN_ADD_1_1_CRY_9,
    O => N_1397);
R1IN_ADD_1_1_CRY_10_Z6416: MUXCY_L port map (
    DI => R1IN_3(42),
    CI => R1IN_ADD_1_1_CRY_9,
    S => R1IN_ADD_1_1_AXB_10,
    LO => R1IN_ADD_1_1_CRY_10);
R1IN_ADD_1_1_S_9: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_9,
    CI => R1IN_ADD_1_1_CRY_8,
    O => N_1395);
R1IN_ADD_1_1_CRY_9_Z6418: MUXCY_L port map (
    DI => R1IN_3(41),
    CI => R1IN_ADD_1_1_CRY_8,
    S => R1IN_ADD_1_1_AXB_9,
    LO => R1IN_ADD_1_1_CRY_9);
R1IN_ADD_1_1_S_8: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_8,
    CI => R1IN_ADD_1_1_CRY_7,
    O => N_1393);
R1IN_ADD_1_1_CRY_8_Z6420: MUXCY_L port map (
    DI => R1IN_3(40),
    CI => R1IN_ADD_1_1_CRY_7,
    S => R1IN_ADD_1_1_AXB_8,
    LO => R1IN_ADD_1_1_CRY_8);
R1IN_ADD_1_1_S_7: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_7,
    CI => R1IN_ADD_1_1_CRY_6,
    O => N_1391);
R1IN_ADD_1_1_CRY_7_Z6422: MUXCY_L port map (
    DI => R1IN_3(39),
    CI => R1IN_ADD_1_1_CRY_6,
    S => R1IN_ADD_1_1_AXB_7,
    LO => R1IN_ADD_1_1_CRY_7);
R1IN_ADD_1_1_S_6: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_6,
    CI => R1IN_ADD_1_1_CRY_5,
    O => N_1389);
R1IN_ADD_1_1_CRY_6_Z6424: MUXCY_L port map (
    DI => R1IN_3(38),
    CI => R1IN_ADD_1_1_CRY_5,
    S => R1IN_ADD_1_1_AXB_6,
    LO => R1IN_ADD_1_1_CRY_6);
R1IN_ADD_1_1_S_5: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_5,
    CI => R1IN_ADD_1_1_CRY_4,
    O => N_1387);
R1IN_ADD_1_1_CRY_5_Z6426: MUXCY_L port map (
    DI => R1IN_3(37),
    CI => R1IN_ADD_1_1_CRY_4,
    S => R1IN_ADD_1_1_AXB_5,
    LO => R1IN_ADD_1_1_CRY_5);
R1IN_ADD_1_1_S_4: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_4,
    CI => R1IN_ADD_1_1_CRY_3,
    O => N_1385);
R1IN_ADD_1_1_CRY_4_Z6428: MUXCY_L port map (
    DI => R1IN_3(36),
    CI => R1IN_ADD_1_1_CRY_3,
    S => R1IN_ADD_1_1_AXB_4,
    LO => R1IN_ADD_1_1_CRY_4);
R1IN_ADD_1_1_S_3: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_3,
    CI => R1IN_ADD_1_1_CRY_2,
    O => N_1383);
R1IN_ADD_1_1_CRY_3_Z6430: MUXCY_L port map (
    DI => R1IN_3(35),
    CI => R1IN_ADD_1_1_CRY_2,
    S => R1IN_ADD_1_1_AXB_3,
    LO => R1IN_ADD_1_1_CRY_3);
R1IN_ADD_1_1_S_2: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_2,
    CI => R1IN_ADD_1_1_CRY_1,
    O => N_1381);
R1IN_ADD_1_1_CRY_2_Z6432: MUXCY_L port map (
    DI => R1IN_3(34),
    CI => R1IN_ADD_1_1_CRY_1,
    S => R1IN_ADD_1_1_AXB_2,
    LO => R1IN_ADD_1_1_CRY_2);
R1IN_ADD_1_1_S_1: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_1,
    CI => R1IN_ADD_1_1_CRY_0,
    O => N_1379);
R1IN_ADD_1_1_CRY_1_Z6434: MUXCY_L port map (
    DI => R1IN_3(33),
    CI => R1IN_ADD_1_1_CRY_0,
    S => R1IN_ADD_1_1_AXB_1,
    LO => R1IN_ADD_1_1_CRY_1);
R1IN_ADD_1_1_CRY_0_Z6435: MUXCY_L port map (
    DI => R1IN_3(32),
    CI => NN_1,
    S => R1IN_ADD_1_1_AXB_0,
    LO => R1IN_ADD_1_1_CRY_0);
R1IN_ADD_1_0_S_31: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_31,
    CI => R1IN_ADD_1_0_CRY_30,
    O => R1IN_ADD_1(31));
R1IN_ADD_1_0_CRY_31_Z6437: MUXCY port map (
    DI => R1IN_3(31),
    CI => R1IN_ADD_1_0_CRY_30,
    S => R1IN_ADD_1_0_AXB_31,
    O => R1IN_ADD_1_0_CRY_31);
R1IN_ADD_1_0_S_30: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_30,
    CI => R1IN_ADD_1_0_CRY_29,
    O => R1IN_ADD_1(30));
R1IN_ADD_1_0_CRY_30_Z6439: MUXCY_L port map (
    DI => R1IN_3(30),
    CI => R1IN_ADD_1_0_CRY_29,
    S => R1IN_ADD_1_0_AXB_30,
    LO => R1IN_ADD_1_0_CRY_30);
R1IN_ADD_1_0_S_29: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_29,
    CI => R1IN_ADD_1_0_CRY_28,
    O => R1IN_ADD_1(29));
R1IN_ADD_1_0_CRY_29_Z6441: MUXCY_L port map (
    DI => R1IN_3(29),
    CI => R1IN_ADD_1_0_CRY_28,
    S => R1IN_ADD_1_0_AXB_29,
    LO => R1IN_ADD_1_0_CRY_29);
R1IN_ADD_1_0_S_28: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_28,
    CI => R1IN_ADD_1_0_CRY_27,
    O => R1IN_ADD_1(28));
R1IN_ADD_1_0_CRY_28_Z6443: MUXCY_L port map (
    DI => R1IN_3(28),
    CI => R1IN_ADD_1_0_CRY_27,
    S => R1IN_ADD_1_0_AXB_28,
    LO => R1IN_ADD_1_0_CRY_28);
R1IN_ADD_1_0_S_27: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_27,
    CI => R1IN_ADD_1_0_CRY_26,
    O => R1IN_ADD_1(27));
R1IN_ADD_1_0_CRY_27_Z6445: MUXCY_L port map (
    DI => R1IN_3(27),
    CI => R1IN_ADD_1_0_CRY_26,
    S => R1IN_ADD_1_0_AXB_27,
    LO => R1IN_ADD_1_0_CRY_27);
R1IN_ADD_1_0_S_26: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_26,
    CI => R1IN_ADD_1_0_CRY_25,
    O => R1IN_ADD_1(26));
R1IN_ADD_1_0_CRY_26_Z6447: MUXCY_L port map (
    DI => R1IN_3(26),
    CI => R1IN_ADD_1_0_CRY_25,
    S => R1IN_ADD_1_0_AXB_26,
    LO => R1IN_ADD_1_0_CRY_26);
R1IN_ADD_1_0_S_25: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_25,
    CI => R1IN_ADD_1_0_CRY_24,
    O => R1IN_ADD_1(25));
R1IN_ADD_1_0_CRY_25_Z6449: MUXCY_L port map (
    DI => R1IN_3(25),
    CI => R1IN_ADD_1_0_CRY_24,
    S => R1IN_ADD_1_0_AXB_25,
    LO => R1IN_ADD_1_0_CRY_25);
R1IN_ADD_1_0_S_24: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_24,
    CI => R1IN_ADD_1_0_CRY_23,
    O => R1IN_ADD_1(24));
R1IN_ADD_1_0_CRY_24_Z6451: MUXCY_L port map (
    DI => R1IN_3(24),
    CI => R1IN_ADD_1_0_CRY_23,
    S => R1IN_ADD_1_0_AXB_24,
    LO => R1IN_ADD_1_0_CRY_24);
R1IN_ADD_1_0_S_23: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_23,
    CI => R1IN_ADD_1_0_CRY_22,
    O => R1IN_ADD_1(23));
R1IN_ADD_1_0_CRY_23_Z6453: MUXCY_L port map (
    DI => R1IN_3(23),
    CI => R1IN_ADD_1_0_CRY_22,
    S => R1IN_ADD_1_0_AXB_23,
    LO => R1IN_ADD_1_0_CRY_23);
R1IN_ADD_1_0_S_22: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_22,
    CI => R1IN_ADD_1_0_CRY_21,
    O => R1IN_ADD_1(22));
R1IN_ADD_1_0_CRY_22_Z6455: MUXCY_L port map (
    DI => R1IN_3(22),
    CI => R1IN_ADD_1_0_CRY_21,
    S => R1IN_ADD_1_0_AXB_22,
    LO => R1IN_ADD_1_0_CRY_22);
R1IN_ADD_1_0_S_21: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_21,
    CI => R1IN_ADD_1_0_CRY_20,
    O => R1IN_ADD_1(21));
R1IN_ADD_1_0_CRY_21_Z6457: MUXCY_L port map (
    DI => R1IN_3(21),
    CI => R1IN_ADD_1_0_CRY_20,
    S => R1IN_ADD_1_0_AXB_21,
    LO => R1IN_ADD_1_0_CRY_21);
R1IN_ADD_1_0_S_20: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_20,
    CI => R1IN_ADD_1_0_CRY_19,
    O => R1IN_ADD_1(20));
R1IN_ADD_1_0_CRY_20_Z6459: MUXCY_L port map (
    DI => R1IN_3(20),
    CI => R1IN_ADD_1_0_CRY_19,
    S => R1IN_ADD_1_0_AXB_20,
    LO => R1IN_ADD_1_0_CRY_20);
R1IN_ADD_1_0_S_19: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_19,
    CI => R1IN_ADD_1_0_CRY_18,
    O => R1IN_ADD_1(19));
R1IN_ADD_1_0_CRY_19_Z6461: MUXCY_L port map (
    DI => R1IN_3(19),
    CI => R1IN_ADD_1_0_CRY_18,
    S => R1IN_ADD_1_0_AXB_19,
    LO => R1IN_ADD_1_0_CRY_19);
R1IN_ADD_1_0_S_18: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_18,
    CI => R1IN_ADD_1_0_CRY_17,
    O => R1IN_ADD_1(18));
R1IN_ADD_1_0_CRY_18_Z6463: MUXCY_L port map (
    DI => R1IN_3(18),
    CI => R1IN_ADD_1_0_CRY_17,
    S => R1IN_ADD_1_0_AXB_18,
    LO => R1IN_ADD_1_0_CRY_18);
R1IN_ADD_1_0_S_17: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_17,
    CI => R1IN_ADD_1_0_CRY_16,
    O => R1IN_ADD_1(17));
R1IN_ADD_1_0_CRY_17_Z6465: MUXCY_L port map (
    DI => R1IN_3(17),
    CI => R1IN_ADD_1_0_CRY_16,
    S => R1IN_ADD_1_0_AXB_17,
    LO => R1IN_ADD_1_0_CRY_17);
R1IN_ADD_1_0_S_16: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_16,
    CI => R1IN_ADD_1_0_CRY_15,
    O => R1IN_ADD_1(16));
R1IN_ADD_1_0_CRY_16_Z6467: MUXCY_L port map (
    DI => R1IN_2F_RETO(16),
    CI => R1IN_ADD_1_0_CRY_15,
    S => R1IN_ADD_1_0_AXB_16,
    LO => R1IN_ADD_1_0_CRY_16);
R1IN_ADD_1_0_S_15: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_15,
    CI => R1IN_ADD_1_0_CRY_14,
    O => R1IN_ADD_1(15));
R1IN_ADD_1_0_CRY_15_Z6469: MUXCY_L port map (
    DI => R1IN_2F_RETO(15),
    CI => R1IN_ADD_1_0_CRY_14,
    S => R1IN_ADD_1_0_AXB_15,
    LO => R1IN_ADD_1_0_CRY_15);
R1IN_ADD_1_0_S_14: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_14,
    CI => R1IN_ADD_1_0_CRY_13,
    O => R1IN_ADD_1(14));
R1IN_ADD_1_0_CRY_14_Z6471: MUXCY_L port map (
    DI => R1IN_2F_RETO(14),
    CI => R1IN_ADD_1_0_CRY_13,
    S => R1IN_ADD_1_0_AXB_14,
    LO => R1IN_ADD_1_0_CRY_14);
R1IN_ADD_1_0_S_13: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_13,
    CI => R1IN_ADD_1_0_CRY_12,
    O => R1IN_ADD_1(13));
R1IN_ADD_1_0_CRY_13_Z6473: MUXCY_L port map (
    DI => R1IN_2F_RETO(13),
    CI => R1IN_ADD_1_0_CRY_12,
    S => R1IN_ADD_1_0_AXB_13,
    LO => R1IN_ADD_1_0_CRY_13);
R1IN_ADD_1_0_S_12: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_12,
    CI => R1IN_ADD_1_0_CRY_11,
    O => R1IN_ADD_1(12));
R1IN_ADD_1_0_CRY_12_Z6475: MUXCY_L port map (
    DI => R1IN_2F_RETO(12),
    CI => R1IN_ADD_1_0_CRY_11,
    S => R1IN_ADD_1_0_AXB_12,
    LO => R1IN_ADD_1_0_CRY_12);
R1IN_ADD_1_0_S_11: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_11,
    CI => R1IN_ADD_1_0_CRY_10,
    O => R1IN_ADD_1(11));
R1IN_ADD_1_0_CRY_11_Z6477: MUXCY_L port map (
    DI => R1IN_2F_RETO(11),
    CI => R1IN_ADD_1_0_CRY_10,
    S => R1IN_ADD_1_0_AXB_11,
    LO => R1IN_ADD_1_0_CRY_11);
R1IN_ADD_1_0_S_10: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_10,
    CI => R1IN_ADD_1_0_CRY_9,
    O => R1IN_ADD_1(10));
R1IN_ADD_1_0_CRY_10_Z6479: MUXCY_L port map (
    DI => R1IN_2F_RETO(10),
    CI => R1IN_ADD_1_0_CRY_9,
    S => R1IN_ADD_1_0_AXB_10,
    LO => R1IN_ADD_1_0_CRY_10);
R1IN_ADD_1_0_S_9: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_9,
    CI => R1IN_ADD_1_0_CRY_8,
    O => R1IN_ADD_1(9));
R1IN_ADD_1_0_CRY_9_Z6481: MUXCY_L port map (
    DI => R1IN_2F_RETO(9),
    CI => R1IN_ADD_1_0_CRY_8,
    S => R1IN_ADD_1_0_AXB_9,
    LO => R1IN_ADD_1_0_CRY_9);
R1IN_ADD_1_0_S_8: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_8,
    CI => R1IN_ADD_1_0_CRY_7,
    O => R1IN_ADD_1(8));
R1IN_ADD_1_0_CRY_8_Z6483: MUXCY_L port map (
    DI => R1IN_2F_RETO(8),
    CI => R1IN_ADD_1_0_CRY_7,
    S => R1IN_ADD_1_0_AXB_8,
    LO => R1IN_ADD_1_0_CRY_8);
R1IN_ADD_1_0_S_7: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_7,
    CI => R1IN_ADD_1_0_CRY_6,
    O => R1IN_ADD_1(7));
R1IN_ADD_1_0_CRY_7_Z6485: MUXCY_L port map (
    DI => R1IN_2F_RETO(7),
    CI => R1IN_ADD_1_0_CRY_6,
    S => R1IN_ADD_1_0_AXB_7,
    LO => R1IN_ADD_1_0_CRY_7);
R1IN_ADD_1_0_S_6: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_6,
    CI => R1IN_ADD_1_0_CRY_5,
    O => R1IN_ADD_1(6));
R1IN_ADD_1_0_CRY_6_Z6487: MUXCY_L port map (
    DI => R1IN_2F_RETO(6),
    CI => R1IN_ADD_1_0_CRY_5,
    S => R1IN_ADD_1_0_AXB_6,
    LO => R1IN_ADD_1_0_CRY_6);
R1IN_ADD_1_0_S_5: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_5,
    CI => R1IN_ADD_1_0_CRY_4,
    O => R1IN_ADD_1(5));
R1IN_ADD_1_0_CRY_5_Z6489: MUXCY_L port map (
    DI => R1IN_2F_RETO(5),
    CI => R1IN_ADD_1_0_CRY_4,
    S => R1IN_ADD_1_0_AXB_5,
    LO => R1IN_ADD_1_0_CRY_5);
R1IN_ADD_1_0_S_4: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_4,
    CI => R1IN_ADD_1_0_CRY_3,
    O => R1IN_ADD_1(4));
R1IN_ADD_1_0_CRY_4_Z6491: MUXCY_L port map (
    DI => R1IN_2F_RETO(4),
    CI => R1IN_ADD_1_0_CRY_3,
    S => R1IN_ADD_1_0_AXB_4,
    LO => R1IN_ADD_1_0_CRY_4);
R1IN_ADD_1_0_S_3: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_3,
    CI => R1IN_ADD_1_0_CRY_2,
    O => R1IN_ADD_1(3));
R1IN_ADD_1_0_CRY_3_Z6493: MUXCY_L port map (
    DI => R1IN_2F_RETO(3),
    CI => R1IN_ADD_1_0_CRY_2,
    S => R1IN_ADD_1_0_AXB_3,
    LO => R1IN_ADD_1_0_CRY_3);
R1IN_ADD_1_0_S_2: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_2,
    CI => R1IN_ADD_1_0_CRY_1,
    O => R1IN_ADD_1(2));
R1IN_ADD_1_0_CRY_2_Z6495: MUXCY_L port map (
    DI => R1IN_2F_RETO(2),
    CI => R1IN_ADD_1_0_CRY_1,
    S => R1IN_ADD_1_0_AXB_2,
    LO => R1IN_ADD_1_0_CRY_2);
R1IN_ADD_1_0_S_1: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_1,
    CI => R1IN_ADD_1_0_CRY_0,
    O => R1IN_ADD_1(1));
R1IN_ADD_1_0_CRY_1_Z6497: MUXCY_L port map (
    DI => R1IN_2F_RETO(1),
    CI => R1IN_ADD_1_0_CRY_0,
    S => R1IN_ADD_1_0_AXB_1,
    LO => R1IN_ADD_1_0_CRY_1);
R1IN_ADD_1_0_CRY_0_Z6498: MUXCY_L port map (
    DI => R1IN_2F_RETO(0),
    CI => NN_1,
    S => R1IN_ADD_1(0),
    LO => R1IN_ADD_1_0_CRY_0);
R1IN_4_ADD_2_1_0_S_34: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_34,
    CI => R1IN_4_ADD_2_1_0_CRY_33,
    O => N_1556);
R1IN_4_ADD_2_1_0_S_33: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_33,
    CI => R1IN_4_ADD_2_1_0_CRY_32,
    O => N_1555);
R1IN_4_ADD_2_1_0_CRY_33_Z6501: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_32,
    S => R1IN_4_ADD_2_1_0_AXB_33,
    LO => R1IN_4_ADD_2_1_0_CRY_33);
R1IN_4_ADD_2_1_0_S_32: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_32,
    CI => R1IN_4_ADD_2_1_0_CRY_31,
    O => N_1554);
R1IN_4_ADD_2_1_0_CRY_32_Z6503: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_31,
    S => R1IN_4_ADD_2_1_0_AXB_32,
    LO => R1IN_4_ADD_2_1_0_CRY_32);
R1IN_4_ADD_2_1_0_S_31: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_31,
    CI => R1IN_4_ADD_2_1_0_CRY_30,
    O => N_1553);
R1IN_4_ADD_2_1_0_CRY_31_Z6505: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_30,
    S => R1IN_4_ADD_2_1_0_AXB_31,
    LO => R1IN_4_ADD_2_1_0_CRY_31);
R1IN_4_ADD_2_1_0_S_30: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_30,
    CI => R1IN_4_ADD_2_1_0_CRY_29,
    O => N_1552);
R1IN_4_ADD_2_1_0_CRY_30_Z6507: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_29,
    S => R1IN_4_ADD_2_1_0_AXB_30,
    LO => R1IN_4_ADD_2_1_0_CRY_30);
R1IN_4_ADD_2_1_0_S_29: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_29,
    CI => R1IN_4_ADD_2_1_0_CRY_28,
    O => N_1551);
R1IN_4_ADD_2_1_0_CRY_29_Z6509: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_28,
    S => R1IN_4_ADD_2_1_0_AXB_29,
    LO => R1IN_4_ADD_2_1_0_CRY_29);
R1IN_4_ADD_2_1_0_S_28: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_28,
    CI => R1IN_4_ADD_2_1_0_CRY_27,
    O => N_1550);
R1IN_4_ADD_2_1_0_CRY_28_Z6511: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_27,
    S => R1IN_4_ADD_2_1_0_AXB_28,
    LO => R1IN_4_ADD_2_1_0_CRY_28);
R1IN_4_ADD_2_1_0_S_27: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_27,
    CI => R1IN_4_ADD_2_1_0_CRY_26,
    O => N_1549);
R1IN_4_ADD_2_1_0_CRY_27_Z6513: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_26,
    S => R1IN_4_ADD_2_1_0_AXB_27,
    LO => R1IN_4_ADD_2_1_0_CRY_27);
R1IN_4_ADD_2_1_0_S_26: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_26,
    CI => R1IN_4_ADD_2_1_0_CRY_25,
    O => N_1548);
R1IN_4_ADD_2_1_0_CRY_26_Z6515: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_25,
    S => R1IN_4_ADD_2_1_0_AXB_26,
    LO => R1IN_4_ADD_2_1_0_CRY_26);
R1IN_4_ADD_2_1_0_S_25: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_25,
    CI => R1IN_4_ADD_2_1_0_CRY_24,
    O => N_1547);
R1IN_4_ADD_2_1_0_CRY_25_Z6517: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_24,
    S => R1IN_4_ADD_2_1_0_AXB_25,
    LO => R1IN_4_ADD_2_1_0_CRY_25);
R1IN_4_ADD_2_1_0_S_24: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_24,
    CI => R1IN_4_ADD_2_1_0_CRY_23,
    O => N_1546);
R1IN_4_ADD_2_1_0_CRY_24_Z6519: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_23,
    S => R1IN_4_ADD_2_1_0_AXB_24,
    LO => R1IN_4_ADD_2_1_0_CRY_24);
R1IN_4_ADD_2_1_0_S_23: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_23,
    CI => R1IN_4_ADD_2_1_0_CRY_22,
    O => N_1545);
R1IN_4_ADD_2_1_0_CRY_23_Z6521: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_22,
    S => R1IN_4_ADD_2_1_0_AXB_23,
    LO => R1IN_4_ADD_2_1_0_CRY_23);
R1IN_4_ADD_2_1_0_S_22: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_22,
    CI => R1IN_4_ADD_2_1_0_CRY_21,
    O => N_1544);
R1IN_4_ADD_2_1_0_CRY_22_Z6523: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_21,
    S => R1IN_4_ADD_2_1_0_AXB_22,
    LO => R1IN_4_ADD_2_1_0_CRY_22);
R1IN_4_ADD_2_1_0_S_21: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_21,
    CI => R1IN_4_ADD_2_1_0_CRY_20,
    O => N_1543);
R1IN_4_ADD_2_1_0_CRY_21_Z6525: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_20,
    S => R1IN_4_ADD_2_1_0_AXB_21,
    LO => R1IN_4_ADD_2_1_0_CRY_21);
R1IN_4_ADD_2_1_0_S_20: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_20,
    CI => R1IN_4_ADD_2_1_0_CRY_19,
    O => N_1542);
R1IN_4_ADD_2_1_0_CRY_20_Z6527: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_19,
    S => R1IN_4_ADD_2_1_0_AXB_20,
    LO => R1IN_4_ADD_2_1_0_CRY_20);
R1IN_4_ADD_2_1_0_S_19: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_19,
    CI => R1IN_4_ADD_2_1_0_CRY_18,
    O => N_1541);
R1IN_4_ADD_2_1_0_CRY_19_Z6529: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_18,
    S => R1IN_4_ADD_2_1_0_AXB_19,
    LO => R1IN_4_ADD_2_1_0_CRY_19);
R1IN_4_ADD_2_1_0_S_18: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_18,
    CI => R1IN_4_ADD_2_1_0_CRY_17,
    O => N_1540);
R1IN_4_ADD_2_1_0_CRY_18_Z6531: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_17,
    S => R1IN_4_ADD_2_1_0_AXB_18,
    LO => R1IN_4_ADD_2_1_0_CRY_18);
R1IN_4_ADD_2_1_0_S_17: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_17,
    CI => R1IN_4_ADD_2_1_0_CRY_16,
    O => N_1539);
R1IN_4_ADD_2_1_0_CRY_17_Z6533: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_16,
    S => R1IN_4_ADD_2_1_0_AXB_17,
    LO => R1IN_4_ADD_2_1_0_CRY_17);
R1IN_4_ADD_2_1_0_S_16: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_16,
    CI => R1IN_4_ADD_2_1_0_CRY_15,
    O => N_1538);
R1IN_4_ADD_2_1_0_CRY_16_Z6535: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_15,
    S => R1IN_4_ADD_2_1_0_AXB_16,
    LO => R1IN_4_ADD_2_1_0_CRY_16);
R1IN_4_ADD_2_1_0_S_15: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_15,
    CI => R1IN_4_ADD_2_1_0_CRY_14,
    O => N_1537);
R1IN_4_ADD_2_1_0_CRY_15_Z6537: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_14,
    S => R1IN_4_ADD_2_1_0_AXB_15,
    LO => R1IN_4_ADD_2_1_0_CRY_15);
R1IN_4_ADD_2_1_0_S_14: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_14,
    CI => R1IN_4_ADD_2_1_0_CRY_13,
    O => N_1536);
R1IN_4_ADD_2_1_0_CRY_14_Z6539: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_13,
    S => R1IN_4_ADD_2_1_0_AXB_14,
    LO => R1IN_4_ADD_2_1_0_CRY_14);
R1IN_4_ADD_2_1_0_S_13: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_13,
    CI => R1IN_4_ADD_2_1_0_CRY_12,
    O => N_1535);
R1IN_4_ADD_2_1_0_CRY_13_Z6541: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_12,
    S => R1IN_4_ADD_2_1_0_AXB_13,
    LO => R1IN_4_ADD_2_1_0_CRY_13);
R1IN_4_ADD_2_1_0_S_12: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_12,
    CI => R1IN_4_ADD_2_1_0_CRY_11,
    O => N_1534);
R1IN_4_ADD_2_1_0_CRY_12_Z6543: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_11,
    S => R1IN_4_ADD_2_1_0_AXB_12,
    LO => R1IN_4_ADD_2_1_0_CRY_12);
R1IN_4_ADD_2_1_0_S_11: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_11,
    CI => R1IN_4_ADD_2_1_0_CRY_10,
    O => N_1533);
R1IN_4_ADD_2_1_0_CRY_11_Z6545: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_10,
    S => R1IN_4_ADD_2_1_0_AXB_11,
    LO => R1IN_4_ADD_2_1_0_CRY_11);
R1IN_4_ADD_2_1_0_S_10: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_10,
    CI => R1IN_4_ADD_2_1_0_CRY_9,
    O => N_1532);
R1IN_4_ADD_2_1_0_CRY_10_Z6547: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_9,
    S => R1IN_4_ADD_2_1_0_AXB_10,
    LO => R1IN_4_ADD_2_1_0_CRY_10);
R1IN_4_ADD_2_1_0_S_9: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_9,
    CI => R1IN_4_ADD_2_1_0_CRY_8,
    O => N_1531);
R1IN_4_ADD_2_1_0_CRY_9_Z6549: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_8,
    S => R1IN_4_ADD_2_1_0_AXB_9,
    LO => R1IN_4_ADD_2_1_0_CRY_9);
R1IN_4_ADD_2_1_0_S_8: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_8,
    CI => R1IN_4_ADD_2_1_0_CRY_7,
    O => N_1530);
R1IN_4_ADD_2_1_0_CRY_8_Z6551: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(44),
    CI => R1IN_4_ADD_2_1_0_CRY_7,
    S => R1IN_4_ADD_2_1_0_AXB_8,
    LO => R1IN_4_ADD_2_1_0_CRY_8);
R1IN_4_ADD_2_1_0_S_7: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_7,
    CI => R1IN_4_ADD_2_1_0_CRY_6,
    O => N_1529);
R1IN_4_ADD_2_1_0_CRY_7_Z6553: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(43),
    CI => R1IN_4_ADD_2_1_0_CRY_6,
    S => R1IN_4_ADD_2_1_0_AXB_7,
    LO => R1IN_4_ADD_2_1_0_CRY_7);
R1IN_4_ADD_2_1_0_S_6: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_6,
    CI => R1IN_4_ADD_2_1_0_CRY_5,
    O => N_1528);
R1IN_4_ADD_2_1_0_CRY_6_Z6555: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(42),
    CI => R1IN_4_ADD_2_1_0_CRY_5,
    S => R1IN_4_ADD_2_1_0_AXB_6,
    LO => R1IN_4_ADD_2_1_0_CRY_6);
R1IN_4_ADD_2_1_0_S_5: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_5,
    CI => R1IN_4_ADD_2_1_0_CRY_4,
    O => N_1527);
R1IN_4_ADD_2_1_0_CRY_5_Z6557: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(41),
    CI => R1IN_4_ADD_2_1_0_CRY_4,
    S => R1IN_4_ADD_2_1_0_AXB_5,
    LO => R1IN_4_ADD_2_1_0_CRY_5);
R1IN_4_ADD_2_1_0_S_4: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_4,
    CI => R1IN_4_ADD_2_1_0_CRY_3,
    O => N_1526);
R1IN_4_ADD_2_1_0_CRY_4_Z6559: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(40),
    CI => R1IN_4_ADD_2_1_0_CRY_3,
    S => R1IN_4_ADD_2_1_0_AXB_4,
    LO => R1IN_4_ADD_2_1_0_CRY_4);
R1IN_4_ADD_2_1_0_S_3: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_3,
    CI => R1IN_4_ADD_2_1_0_CRY_2,
    O => N_1525);
R1IN_4_ADD_2_1_0_CRY_3_Z6561: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(39),
    CI => R1IN_4_ADD_2_1_0_CRY_2,
    S => R1IN_4_ADD_2_1_0_AXB_3,
    LO => R1IN_4_ADD_2_1_0_CRY_3);
R1IN_4_ADD_2_1_0_S_2: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_2,
    CI => R1IN_4_ADD_2_1_0_CRY_1,
    O => N_1524);
R1IN_4_ADD_2_1_0_CRY_2_Z6563: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(38),
    CI => R1IN_4_ADD_2_1_0_CRY_1,
    S => R1IN_4_ADD_2_1_0_AXB_2,
    LO => R1IN_4_ADD_2_1_0_CRY_2);
R1IN_4_ADD_2_1_0_S_1: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_1,
    CI => R1IN_4_ADD_2_1_0_CRY_0,
    O => N_1523);
R1IN_4_ADD_2_1_0_CRY_1_Z6565: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(37),
    CI => R1IN_4_ADD_2_1_0_CRY_0,
    S => R1IN_4_ADD_2_1_0_AXB_1,
    LO => R1IN_4_ADD_2_1_0_CRY_1);
R1IN_4_ADD_2_1_0_CRY_0_Z6566: MUXCY_L port map (
    DI => R1IN_4_ADD_2_1_RETO,
    CI => NN_2,
    S => R1IN_4_ADD_2_1_0_AXB_0,
    LO => R1IN_4_ADD_2_1_0_CRY_0);
R1IN_4_ADD_2_1_S_34: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_34,
    CI => R1IN_4_ADD_2_1_CRY_33,
    O => N_1511);
R1IN_4_ADD_2_1_S_33: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_33,
    CI => R1IN_4_ADD_2_1_CRY_32,
    O => N_1509);
R1IN_4_ADD_2_1_CRY_33_Z6569: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_32,
    S => R1IN_4_ADD_2_1_AXB_33,
    LO => R1IN_4_ADD_2_1_CRY_33);
R1IN_4_ADD_2_1_S_32: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_32,
    CI => R1IN_4_ADD_2_1_CRY_31,
    O => N_1507);
R1IN_4_ADD_2_1_CRY_32_Z6571: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_31,
    S => R1IN_4_ADD_2_1_AXB_32,
    LO => R1IN_4_ADD_2_1_CRY_32);
R1IN_4_ADD_2_1_S_31: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_31,
    CI => R1IN_4_ADD_2_1_CRY_30,
    O => N_1505);
R1IN_4_ADD_2_1_CRY_31_Z6573: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_30,
    S => R1IN_4_ADD_2_1_AXB_31,
    LO => R1IN_4_ADD_2_1_CRY_31);
R1IN_4_ADD_2_1_S_30: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_30,
    CI => R1IN_4_ADD_2_1_CRY_29,
    O => N_1503);
R1IN_4_ADD_2_1_CRY_30_Z6575: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_29,
    S => R1IN_4_ADD_2_1_AXB_30,
    LO => R1IN_4_ADD_2_1_CRY_30);
R1IN_4_ADD_2_1_S_29: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_29,
    CI => R1IN_4_ADD_2_1_CRY_28,
    O => N_1501);
R1IN_4_ADD_2_1_CRY_29_Z6577: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_28,
    S => R1IN_4_ADD_2_1_AXB_29,
    LO => R1IN_4_ADD_2_1_CRY_29);
R1IN_4_ADD_2_1_S_28: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_28,
    CI => R1IN_4_ADD_2_1_CRY_27,
    O => N_1499);
R1IN_4_ADD_2_1_CRY_28_Z6579: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_27,
    S => R1IN_4_ADD_2_1_AXB_28,
    LO => R1IN_4_ADD_2_1_CRY_28);
R1IN_4_ADD_2_1_S_27: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_27,
    CI => R1IN_4_ADD_2_1_CRY_26,
    O => N_1497);
R1IN_4_ADD_2_1_CRY_27_Z6581: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_26,
    S => R1IN_4_ADD_2_1_AXB_27,
    LO => R1IN_4_ADD_2_1_CRY_27);
R1IN_4_ADD_2_1_S_26: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_26,
    CI => R1IN_4_ADD_2_1_CRY_25,
    O => N_1495);
R1IN_4_ADD_2_1_CRY_26_Z6583: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_25,
    S => R1IN_4_ADD_2_1_AXB_26,
    LO => R1IN_4_ADD_2_1_CRY_26);
R1IN_4_ADD_2_1_S_25: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_25,
    CI => R1IN_4_ADD_2_1_CRY_24,
    O => N_1493);
R1IN_4_ADD_2_1_CRY_25_Z6585: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_24,
    S => R1IN_4_ADD_2_1_AXB_25,
    LO => R1IN_4_ADD_2_1_CRY_25);
R1IN_4_ADD_2_1_S_24: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_24,
    CI => R1IN_4_ADD_2_1_CRY_23,
    O => N_1491);
R1IN_4_ADD_2_1_CRY_24_Z6587: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_23,
    S => R1IN_4_ADD_2_1_AXB_24,
    LO => R1IN_4_ADD_2_1_CRY_24);
R1IN_4_ADD_2_1_S_23: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_23,
    CI => R1IN_4_ADD_2_1_CRY_22,
    O => N_1489);
R1IN_4_ADD_2_1_CRY_23_Z6589: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_22,
    S => R1IN_4_ADD_2_1_AXB_23,
    LO => R1IN_4_ADD_2_1_CRY_23);
R1IN_4_ADD_2_1_S_22: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_22,
    CI => R1IN_4_ADD_2_1_CRY_21,
    O => N_1487);
R1IN_4_ADD_2_1_CRY_22_Z6591: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_21,
    S => R1IN_4_ADD_2_1_AXB_22,
    LO => R1IN_4_ADD_2_1_CRY_22);
R1IN_4_ADD_2_1_S_21: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_21,
    CI => R1IN_4_ADD_2_1_CRY_20,
    O => N_1485);
R1IN_4_ADD_2_1_CRY_21_Z6593: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_20,
    S => R1IN_4_ADD_2_1_AXB_21,
    LO => R1IN_4_ADD_2_1_CRY_21);
R1IN_4_ADD_2_1_S_20: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_20,
    CI => R1IN_4_ADD_2_1_CRY_19,
    O => N_1483);
R1IN_4_ADD_2_1_CRY_20_Z6595: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_19,
    S => R1IN_4_ADD_2_1_AXB_20,
    LO => R1IN_4_ADD_2_1_CRY_20);
R1IN_4_ADD_2_1_S_19: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_19,
    CI => R1IN_4_ADD_2_1_CRY_18,
    O => N_1481);
R1IN_4_ADD_2_1_CRY_19_Z6597: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_18,
    S => R1IN_4_ADD_2_1_AXB_19,
    LO => R1IN_4_ADD_2_1_CRY_19);
R1IN_4_ADD_2_1_S_18: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_18,
    CI => R1IN_4_ADD_2_1_CRY_17,
    O => N_1479);
R1IN_4_ADD_2_1_CRY_18_Z6599: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_17,
    S => R1IN_4_ADD_2_1_AXB_18,
    LO => R1IN_4_ADD_2_1_CRY_18);
R1IN_4_ADD_2_1_S_17: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_17,
    CI => R1IN_4_ADD_2_1_CRY_16,
    O => N_1477);
R1IN_4_ADD_2_1_CRY_17_Z6601: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_16,
    S => R1IN_4_ADD_2_1_AXB_17,
    LO => R1IN_4_ADD_2_1_CRY_17);
R1IN_4_ADD_2_1_S_16: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_16,
    CI => R1IN_4_ADD_2_1_CRY_15,
    O => N_1475);
R1IN_4_ADD_2_1_CRY_16_Z6603: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_15,
    S => R1IN_4_ADD_2_1_AXB_16,
    LO => R1IN_4_ADD_2_1_CRY_16);
R1IN_4_ADD_2_1_S_15: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_15,
    CI => R1IN_4_ADD_2_1_CRY_14,
    O => N_1473);
R1IN_4_ADD_2_1_CRY_15_Z6605: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_14,
    S => R1IN_4_ADD_2_1_AXB_15,
    LO => R1IN_4_ADD_2_1_CRY_15);
R1IN_4_ADD_2_1_S_14: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_14,
    CI => R1IN_4_ADD_2_1_CRY_13,
    O => N_1471);
R1IN_4_ADD_2_1_CRY_14_Z6607: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_13,
    S => R1IN_4_ADD_2_1_AXB_14,
    LO => R1IN_4_ADD_2_1_CRY_14);
R1IN_4_ADD_2_1_S_13: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_13,
    CI => R1IN_4_ADD_2_1_CRY_12,
    O => N_1469);
R1IN_4_ADD_2_1_CRY_13_Z6609: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_12,
    S => R1IN_4_ADD_2_1_AXB_13,
    LO => R1IN_4_ADD_2_1_CRY_13);
R1IN_4_ADD_2_1_S_12: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_12,
    CI => R1IN_4_ADD_2_1_CRY_11,
    O => N_1467);
R1IN_4_ADD_2_1_CRY_12_Z6611: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_11,
    S => R1IN_4_ADD_2_1_AXB_12,
    LO => R1IN_4_ADD_2_1_CRY_12);
R1IN_4_ADD_2_1_S_11: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_11,
    CI => R1IN_4_ADD_2_1_CRY_10,
    O => N_1465);
R1IN_4_ADD_2_1_CRY_11_Z6613: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_10,
    S => R1IN_4_ADD_2_1_AXB_11,
    LO => R1IN_4_ADD_2_1_CRY_11);
R1IN_4_ADD_2_1_S_10: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_10,
    CI => R1IN_4_ADD_2_1_CRY_9,
    O => N_1463);
R1IN_4_ADD_2_1_CRY_10_Z6615: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_9,
    S => R1IN_4_ADD_2_1_AXB_10,
    LO => R1IN_4_ADD_2_1_CRY_10);
R1IN_4_ADD_2_1_S_9: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_9,
    CI => R1IN_4_ADD_2_1_CRY_8,
    O => N_1461);
R1IN_4_ADD_2_1_CRY_9_Z6617: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_8,
    S => R1IN_4_ADD_2_1_AXB_9,
    LO => R1IN_4_ADD_2_1_CRY_9);
R1IN_4_ADD_2_1_S_8: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_8,
    CI => R1IN_4_ADD_2_1_CRY_7,
    O => N_1459);
R1IN_4_ADD_2_1_CRY_8_Z6619: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(44),
    CI => R1IN_4_ADD_2_1_CRY_7,
    S => R1IN_4_ADD_2_1_AXB_8,
    LO => R1IN_4_ADD_2_1_CRY_8);
R1IN_4_ADD_2_1_S_7: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_7,
    CI => R1IN_4_ADD_2_1_CRY_6,
    O => N_1457);
R1IN_4_ADD_2_1_CRY_7_Z6621: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(43),
    CI => R1IN_4_ADD_2_1_CRY_6,
    S => R1IN_4_ADD_2_1_AXB_7,
    LO => R1IN_4_ADD_2_1_CRY_7);
R1IN_4_ADD_2_1_S_6: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_6,
    CI => R1IN_4_ADD_2_1_CRY_5,
    O => N_1455);
R1IN_4_ADD_2_1_CRY_6_Z6623: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(42),
    CI => R1IN_4_ADD_2_1_CRY_5,
    S => R1IN_4_ADD_2_1_AXB_6,
    LO => R1IN_4_ADD_2_1_CRY_6);
R1IN_4_ADD_2_1_S_5: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_5,
    CI => R1IN_4_ADD_2_1_CRY_4,
    O => N_1453);
R1IN_4_ADD_2_1_CRY_5_Z6625: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(41),
    CI => R1IN_4_ADD_2_1_CRY_4,
    S => R1IN_4_ADD_2_1_AXB_5,
    LO => R1IN_4_ADD_2_1_CRY_5);
R1IN_4_ADD_2_1_S_4: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_4,
    CI => R1IN_4_ADD_2_1_CRY_3,
    O => N_1451);
R1IN_4_ADD_2_1_CRY_4_Z6627: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(40),
    CI => R1IN_4_ADD_2_1_CRY_3,
    S => R1IN_4_ADD_2_1_AXB_4,
    LO => R1IN_4_ADD_2_1_CRY_4);
R1IN_4_ADD_2_1_S_3: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_3,
    CI => R1IN_4_ADD_2_1_CRY_2,
    O => N_1449);
R1IN_4_ADD_2_1_CRY_3_Z6629: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(39),
    CI => R1IN_4_ADD_2_1_CRY_2,
    S => R1IN_4_ADD_2_1_AXB_3,
    LO => R1IN_4_ADD_2_1_CRY_3);
R1IN_4_ADD_2_1_S_2: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_2,
    CI => R1IN_4_ADD_2_1_CRY_1,
    O => N_1447);
R1IN_4_ADD_2_1_CRY_2_Z6631: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(38),
    CI => R1IN_4_ADD_2_1_CRY_1,
    S => R1IN_4_ADD_2_1_AXB_2,
    LO => R1IN_4_ADD_2_1_CRY_2);
R1IN_4_ADD_2_1_S_1: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_1,
    CI => R1IN_4_ADD_2_1_CRY_0,
    O => N_1445);
R1IN_4_ADD_2_1_CRY_1_Z6633: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(37),
    CI => R1IN_4_ADD_2_1_CRY_0,
    S => R1IN_4_ADD_2_1_AXB_1,
    LO => R1IN_4_ADD_2_1_CRY_1);
R1IN_4_ADD_2_1_CRY_0_Z6634: MUXCY_L port map (
    DI => R1IN_4_ADD_2_1_RETO,
    CI => NN_1,
    S => R1IN_4_ADD_2_1_AXB_0,
    LO => R1IN_4_ADD_2_1_CRY_0);
R1IN_4_ADD_2_0_S_35: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_35,
    CI => R1IN_4_ADD_2_0_CRY_34,
    O => R1IN_4(52));
R1IN_4_ADD_2_0_CRY_35_Z6636: MUXCY port map (
    DI => R1IN_4_ADD_1_RETO(35),
    CI => R1IN_4_ADD_2_0_CRY_34,
    S => R1IN_4_ADD_2_0_AXB_35,
    O => R1IN_4_ADD_2_0_CRY_35);
R1IN_4_ADD_2_0_S_34: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_34,
    CI => R1IN_4_ADD_2_0_CRY_33,
    O => R1IN_4(51));
R1IN_4_ADD_2_0_CRY_34_Z6638: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(34),
    CI => R1IN_4_ADD_2_0_CRY_33,
    S => R1IN_4_ADD_2_0_AXB_34,
    LO => R1IN_4_ADD_2_0_CRY_34);
R1IN_4_ADD_2_0_S_33: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_33,
    CI => R1IN_4_ADD_2_0_CRY_32,
    O => R1IN_4(50));
R1IN_4_ADD_2_0_CRY_33_Z6640: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(33),
    CI => R1IN_4_ADD_2_0_CRY_32,
    S => R1IN_4_ADD_2_0_AXB_33,
    LO => R1IN_4_ADD_2_0_CRY_33);
R1IN_4_ADD_2_0_S_32: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_32,
    CI => R1IN_4_ADD_2_0_CRY_31,
    O => R1IN_4(49));
R1IN_4_ADD_2_0_CRY_32_Z6642: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(32),
    CI => R1IN_4_ADD_2_0_CRY_31,
    S => R1IN_4_ADD_2_0_AXB_32,
    LO => R1IN_4_ADD_2_0_CRY_32);
R1IN_4_ADD_2_0_S_31: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_31,
    CI => R1IN_4_ADD_2_0_CRY_30,
    O => R1IN_4(48));
R1IN_4_ADD_2_0_CRY_31_Z6644: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(31),
    CI => R1IN_4_ADD_2_0_CRY_30,
    S => R1IN_4_ADD_2_0_AXB_31,
    LO => R1IN_4_ADD_2_0_CRY_31);
R1IN_4_ADD_2_0_S_30: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_30,
    CI => R1IN_4_ADD_2_0_CRY_29,
    O => R1IN_4(47));
R1IN_4_ADD_2_0_CRY_30_Z6646: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(30),
    CI => R1IN_4_ADD_2_0_CRY_29,
    S => R1IN_4_ADD_2_0_AXB_30,
    LO => R1IN_4_ADD_2_0_CRY_30);
R1IN_4_ADD_2_0_S_29: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_29,
    CI => R1IN_4_ADD_2_0_CRY_28,
    O => R1IN_4(46));
R1IN_4_ADD_2_0_CRY_29_Z6648: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(29),
    CI => R1IN_4_ADD_2_0_CRY_28,
    S => R1IN_4_ADD_2_0_AXB_29,
    LO => R1IN_4_ADD_2_0_CRY_29);
R1IN_4_ADD_2_0_S_28: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_28,
    CI => R1IN_4_ADD_2_0_CRY_27,
    O => R1IN_4(45));
R1IN_4_ADD_2_0_CRY_28_Z6650: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(28),
    CI => R1IN_4_ADD_2_0_CRY_27,
    S => R1IN_4_ADD_2_0_AXB_28,
    LO => R1IN_4_ADD_2_0_CRY_28);
R1IN_4_ADD_2_0_S_27: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_27,
    CI => R1IN_4_ADD_2_0_CRY_26,
    O => R1IN_4(44));
R1IN_4_ADD_2_0_CRY_27_Z6652: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(27),
    CI => R1IN_4_ADD_2_0_CRY_26,
    S => R1IN_4_ADD_2_0_AXB_27,
    LO => R1IN_4_ADD_2_0_CRY_27);
R1IN_4_ADD_2_0_S_26: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_26,
    CI => R1IN_4_ADD_2_0_CRY_25,
    O => R1IN_4(43));
R1IN_4_ADD_2_0_CRY_26_Z6654: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(26),
    CI => R1IN_4_ADD_2_0_CRY_25,
    S => R1IN_4_ADD_2_0_AXB_26,
    LO => R1IN_4_ADD_2_0_CRY_26);
R1IN_4_ADD_2_0_S_25: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_25,
    CI => R1IN_4_ADD_2_0_CRY_24,
    O => R1IN_4(42));
R1IN_4_ADD_2_0_CRY_25_Z6656: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(25),
    CI => R1IN_4_ADD_2_0_CRY_24,
    S => R1IN_4_ADD_2_0_AXB_25,
    LO => R1IN_4_ADD_2_0_CRY_25);
R1IN_4_ADD_2_0_S_24: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_24,
    CI => R1IN_4_ADD_2_0_CRY_23,
    O => R1IN_4(41));
R1IN_4_ADD_2_0_CRY_24_Z6658: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(24),
    CI => R1IN_4_ADD_2_0_CRY_23,
    S => R1IN_4_ADD_2_0_AXB_24,
    LO => R1IN_4_ADD_2_0_CRY_24);
R1IN_4_ADD_2_0_S_23: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_23,
    CI => R1IN_4_ADD_2_0_CRY_22,
    O => R1IN_4(40));
R1IN_4_ADD_2_0_CRY_23_Z6660: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(23),
    CI => R1IN_4_ADD_2_0_CRY_22,
    S => R1IN_4_ADD_2_0_AXB_23,
    LO => R1IN_4_ADD_2_0_CRY_23);
R1IN_4_ADD_2_0_S_22: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_22,
    CI => R1IN_4_ADD_2_0_CRY_21,
    O => R1IN_4(39));
R1IN_4_ADD_2_0_CRY_22_Z6662: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(22),
    CI => R1IN_4_ADD_2_0_CRY_21,
    S => R1IN_4_ADD_2_0_AXB_22,
    LO => R1IN_4_ADD_2_0_CRY_22);
R1IN_4_ADD_2_0_S_21: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_21,
    CI => R1IN_4_ADD_2_0_CRY_20,
    O => R1IN_4(38));
R1IN_4_ADD_2_0_CRY_21_Z6664: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(21),
    CI => R1IN_4_ADD_2_0_CRY_20,
    S => R1IN_4_ADD_2_0_AXB_21,
    LO => R1IN_4_ADD_2_0_CRY_21);
R1IN_4_ADD_2_0_S_20: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_20,
    CI => R1IN_4_ADD_2_0_CRY_19,
    O => R1IN_4(37));
R1IN_4_ADD_2_0_CRY_20_Z6666: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(20),
    CI => R1IN_4_ADD_2_0_CRY_19,
    S => R1IN_4_ADD_2_0_AXB_20,
    LO => R1IN_4_ADD_2_0_CRY_20);
R1IN_4_ADD_2_0_S_19: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_19,
    CI => R1IN_4_ADD_2_0_CRY_18,
    O => R1IN_4(36));
R1IN_4_ADD_2_0_CRY_19_Z6668: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(19),
    CI => R1IN_4_ADD_2_0_CRY_18,
    S => R1IN_4_ADD_2_0_AXB_19,
    LO => R1IN_4_ADD_2_0_CRY_19);
R1IN_4_ADD_2_0_S_18: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_18,
    CI => R1IN_4_ADD_2_0_CRY_17,
    O => R1IN_4(35));
R1IN_4_ADD_2_0_CRY_18_Z6670: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(18),
    CI => R1IN_4_ADD_2_0_CRY_17,
    S => R1IN_4_ADD_2_0_AXB_18,
    LO => R1IN_4_ADD_2_0_CRY_18);
R1IN_4_ADD_2_0_S_17: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_17,
    CI => R1IN_4_ADD_2_0_CRY_16,
    O => R1IN_4(34));
R1IN_4_ADD_2_0_CRY_17_Z6672: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(17),
    CI => R1IN_4_ADD_2_0_CRY_16,
    S => R1IN_4_ADD_2_0_AXB_17,
    LO => R1IN_4_ADD_2_0_CRY_17);
R1IN_4_ADD_2_0_S_16: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_16,
    CI => R1IN_4_ADD_2_0_CRY_15,
    O => R1IN_4(33));
R1IN_4_ADD_2_0_CRY_16_Z6674: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(16),
    CI => R1IN_4_ADD_2_0_CRY_15,
    S => R1IN_4_ADD_2_0_AXB_16,
    LO => R1IN_4_ADD_2_0_CRY_16);
R1IN_4_ADD_2_0_S_15: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_15,
    CI => R1IN_4_ADD_2_0_CRY_14,
    O => R1IN_4(32));
R1IN_4_ADD_2_0_CRY_15_Z6676: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(15),
    CI => R1IN_4_ADD_2_0_CRY_14,
    S => R1IN_4_ADD_2_0_AXB_15,
    LO => R1IN_4_ADD_2_0_CRY_15);
R1IN_4_ADD_2_0_S_14: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_14,
    CI => R1IN_4_ADD_2_0_CRY_13,
    O => R1IN_4(31));
R1IN_4_ADD_2_0_CRY_14_Z6678: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(14),
    CI => R1IN_4_ADD_2_0_CRY_13,
    S => R1IN_4_ADD_2_0_AXB_14,
    LO => R1IN_4_ADD_2_0_CRY_14);
R1IN_4_ADD_2_0_S_13: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_13,
    CI => R1IN_4_ADD_2_0_CRY_12,
    O => R1IN_4(30));
R1IN_4_ADD_2_0_CRY_13_Z6680: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(13),
    CI => R1IN_4_ADD_2_0_CRY_12,
    S => R1IN_4_ADD_2_0_AXB_13,
    LO => R1IN_4_ADD_2_0_CRY_13);
R1IN_4_ADD_2_0_S_12: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_12,
    CI => R1IN_4_ADD_2_0_CRY_11,
    O => R1IN_4(29));
R1IN_4_ADD_2_0_CRY_12_Z6682: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(12),
    CI => R1IN_4_ADD_2_0_CRY_11,
    S => R1IN_4_ADD_2_0_AXB_12,
    LO => R1IN_4_ADD_2_0_CRY_12);
R1IN_4_ADD_2_0_S_11: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_11,
    CI => R1IN_4_ADD_2_0_CRY_10,
    O => R1IN_4(28));
R1IN_4_ADD_2_0_CRY_11_Z6684: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(11),
    CI => R1IN_4_ADD_2_0_CRY_10,
    S => R1IN_4_ADD_2_0_AXB_11,
    LO => R1IN_4_ADD_2_0_CRY_11);
R1IN_4_ADD_2_0_S_10: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_10,
    CI => R1IN_4_ADD_2_0_CRY_9,
    O => R1IN_4(27));
R1IN_4_ADD_2_0_CRY_10_Z6686: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(10),
    CI => R1IN_4_ADD_2_0_CRY_9,
    S => R1IN_4_ADD_2_0_AXB_10,
    LO => R1IN_4_ADD_2_0_CRY_10);
R1IN_4_ADD_2_0_S_9: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_9,
    CI => R1IN_4_ADD_2_0_CRY_8,
    O => R1IN_4(26));
R1IN_4_ADD_2_0_CRY_9_Z6688: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(9),
    CI => R1IN_4_ADD_2_0_CRY_8,
    S => R1IN_4_ADD_2_0_AXB_9,
    LO => R1IN_4_ADD_2_0_CRY_9);
R1IN_4_ADD_2_0_S_8: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_8,
    CI => R1IN_4_ADD_2_0_CRY_7,
    O => R1IN_4(25));
R1IN_4_ADD_2_0_CRY_8_Z6690: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(8),
    CI => R1IN_4_ADD_2_0_CRY_7,
    S => R1IN_4_ADD_2_0_AXB_8,
    LO => R1IN_4_ADD_2_0_CRY_8);
R1IN_4_ADD_2_0_S_7: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_7,
    CI => R1IN_4_ADD_2_0_CRY_6,
    O => R1IN_4(24));
R1IN_4_ADD_2_0_CRY_7_Z6692: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(7),
    CI => R1IN_4_ADD_2_0_CRY_6,
    S => R1IN_4_ADD_2_0_AXB_7,
    LO => R1IN_4_ADD_2_0_CRY_7);
R1IN_4_ADD_2_0_S_6: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_6,
    CI => R1IN_4_ADD_2_0_CRY_5,
    O => R1IN_4(23));
R1IN_4_ADD_2_0_CRY_6_Z6694: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(6),
    CI => R1IN_4_ADD_2_0_CRY_5,
    S => R1IN_4_ADD_2_0_AXB_6,
    LO => R1IN_4_ADD_2_0_CRY_6);
R1IN_4_ADD_2_0_S_5: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_5,
    CI => R1IN_4_ADD_2_0_CRY_4,
    O => R1IN_4(22));
R1IN_4_ADD_2_0_CRY_5_Z6696: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(5),
    CI => R1IN_4_ADD_2_0_CRY_4,
    S => R1IN_4_ADD_2_0_AXB_5,
    LO => R1IN_4_ADD_2_0_CRY_5);
R1IN_4_ADD_2_0_S_4: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_4,
    CI => R1IN_4_ADD_2_0_CRY_3,
    O => R1IN_4(21));
R1IN_4_ADD_2_0_CRY_4_Z6698: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(4),
    CI => R1IN_4_ADD_2_0_CRY_3,
    S => R1IN_4_ADD_2_0_AXB_4,
    LO => R1IN_4_ADD_2_0_CRY_4);
R1IN_4_ADD_2_0_S_3: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_3,
    CI => R1IN_4_ADD_2_0_CRY_2,
    O => R1IN_4(20));
R1IN_4_ADD_2_0_CRY_3_Z6700: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(3),
    CI => R1IN_4_ADD_2_0_CRY_2,
    S => R1IN_4_ADD_2_0_AXB_3,
    LO => R1IN_4_ADD_2_0_CRY_3);
R1IN_4_ADD_2_0_S_2: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_2,
    CI => R1IN_4_ADD_2_0_CRY_1,
    O => R1IN_4(19));
R1IN_4_ADD_2_0_CRY_2_Z6702: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(2),
    CI => R1IN_4_ADD_2_0_CRY_1,
    S => R1IN_4_ADD_2_0_AXB_2,
    LO => R1IN_4_ADD_2_0_CRY_2);
R1IN_4_ADD_2_0_S_1: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_1,
    CI => R1IN_4_ADD_2_0_CRY_0,
    O => R1IN_4(18));
R1IN_4_ADD_2_0_CRY_1_Z6704: MUXCY_L port map (
    DI => R1IN_4_ADD_1_RETO(1),
    CI => R1IN_4_ADD_2_0_CRY_0,
    S => R1IN_4_ADD_2_0_AXB_1,
    LO => R1IN_4_ADD_2_0_CRY_1);
R1IN_4_ADD_2_0_CRY_0_Z6705: MUXCY_L port map (
    DI => R1IN_4_ADD_2_0_RETO,
    CI => NN_1,
    S => R1IN_4(17),
    LO => R1IN_4_ADD_2_0_CRY_0);
R1IN_4_4_4q190w: DSP48 
generic map(
  AREG => 1,
  BREG => 1,
  CREG => 0,
  PREG => 1,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => A(51),
  A(1) => A(52),
  A(2) => A(53),
  A(3) => A(54),
  A(4) => A(55),
  A(5) => A(56),
  A(6) => A(57),
  A(7) => A(58),
  A(8) => A(59),
  A(9) => A(60),
  A(10) => NN_1,
  A(11) => NN_1,
  A(12) => NN_1,
  A(13) => NN_1,
  A(14) => NN_1,
  A(15) => NN_1,
  A(16) => NN_1,
  A(17) => NN_1,
  B(0) => B(51),
  B(1) => B(52),
  B(2) => B(53),
  B(3) => B(54),
  B(4) => B(55),
  B(5) => B(56),
  B(6) => B(57),
  B(7) => B(58),
  B(8) => B(59),
  B(9) => B(60),
  B(10) => NN_1,
  B(11) => NN_1,
  B(12) => NN_1,
  B(13) => NN_1,
  B(14) => NN_1,
  B(15) => NN_1,
  B(16) => NN_1,
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => NN_1,
  PCIN(1) => NN_1,
  PCIN(2) => NN_1,
  PCIN(3) => NN_1,
  PCIN(4) => NN_1,
  PCIN(5) => NN_1,
  PCIN(6) => NN_1,
  PCIN(7) => NN_1,
  PCIN(8) => NN_1,
  PCIN(9) => NN_1,
  PCIN(10) => NN_1,
  PCIN(11) => NN_1,
  PCIN(12) => NN_1,
  PCIN(13) => NN_1,
  PCIN(14) => NN_1,
  PCIN(15) => NN_1,
  PCIN(16) => NN_1,
  PCIN(17) => NN_1,
  PCIN(18) => NN_1,
  PCIN(19) => NN_1,
  PCIN(20) => NN_1,
  PCIN(21) => NN_1,
  PCIN(22) => NN_1,
  PCIN(23) => NN_1,
  PCIN(24) => NN_1,
  PCIN(25) => NN_1,
  PCIN(26) => NN_1,
  PCIN(27) => NN_1,
  PCIN(28) => NN_1,
  PCIN(29) => NN_1,
  PCIN(30) => NN_1,
  PCIN(31) => NN_1,
  PCIN(32) => NN_1,
  PCIN(33) => NN_1,
  PCIN(34) => NN_1,
  PCIN(35) => NN_1,
  PCIN(36) => NN_1,
  PCIN(37) => NN_1,
  PCIN(38) => NN_1,
  PCIN(39) => NN_1,
  PCIN(40) => NN_1,
  PCIN(41) => NN_1,
  PCIN(42) => NN_1,
  PCIN(43) => NN_1,
  PCIN(44) => NN_1,
  PCIN(45) => NN_1,
  PCIN(46) => NN_1,
  PCIN(47) => NN_1,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_1,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => CLK,
  CEA => EN,
  CEB => EN,
  CEC => NN_1,
  CEP => EN,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_4_4_4_BCOUT(0),
  BCOUT(1) => R1IN_4_4_4_BCOUT(1),
  BCOUT(2) => R1IN_4_4_4_BCOUT(2),
  BCOUT(3) => R1IN_4_4_4_BCOUT(3),
  BCOUT(4) => R1IN_4_4_4_BCOUT(4),
  BCOUT(5) => R1IN_4_4_4_BCOUT(5),
  BCOUT(6) => R1IN_4_4_4_BCOUT(6),
  BCOUT(7) => R1IN_4_4_4_BCOUT(7),
  BCOUT(8) => R1IN_4_4_4_BCOUT(8),
  BCOUT(9) => R1IN_4_4_4_BCOUT(9),
  BCOUT(10) => R1IN_4_4_4_BCOUT(10),
  BCOUT(11) => R1IN_4_4_4_BCOUT(11),
  BCOUT(12) => R1IN_4_4_4_BCOUT(12),
  BCOUT(13) => R1IN_4_4_4_BCOUT(13),
  BCOUT(14) => R1IN_4_4_4_BCOUT(14),
  BCOUT(15) => R1IN_4_4_4_BCOUT(15),
  BCOUT(16) => R1IN_4_4_4_BCOUT(16),
  BCOUT(17) => R1IN_4_4_4_BCOUT(17),
  P(0) => R1IN_4_4_4F_RETO(0),
  P(1) => R1IN_4_4_4F_RETO(1),
  P(2) => R1IN_4_4_4F_RETO(2),
  P(3) => R1IN_4_4_4F_RETO(3),
  P(4) => R1IN_4_4_4F_RETO(4),
  P(5) => R1IN_4_4_4F_RETO(5),
  P(6) => R1IN_4_4_4F_RETO(6),
  P(7) => R1IN_4_4_4F_RETO(7),
  P(8) => R1IN_4_4_4F_RETO(8),
  P(9) => R1IN_4_4_4F_RETO(9),
  P(10) => R1IN_4_4_4F_RETO(10),
  P(11) => R1IN_4_4_4F_RETO(11),
  P(12) => R1IN_4_4_4F_RETO(12),
  P(13) => R1IN_4_4_4F_RETO(13),
  P(14) => R1IN_4_4_4F_RETO(14),
  P(15) => R1IN_4_4_4F_RETO(15),
  P(16) => R1IN_4_4_4F_RETO(16),
  P(17) => R1IN_4_4_4F_RETO(17),
  P(18) => R1IN_4_4_4F_RETO(18),
  P(19) => R1IN_4_4_4F_RETO(19),
  P(20) => R1IN_4_4_4_P(20),
  P(21) => R1IN_4_4_4_P(21),
  P(22) => R1IN_4_4_4_P(22),
  P(23) => R1IN_4_4_4_P(23),
  P(24) => R1IN_4_4_4_P(24),
  P(25) => R1IN_4_4_4_P(25),
  P(26) => R1IN_4_4_4_P(26),
  P(27) => R1IN_4_4_4_P(27),
  P(28) => R1IN_4_4_4_P(28),
  P(29) => R1IN_4_4_4_P(29),
  P(30) => R1IN_4_4_4_P(30),
  P(31) => R1IN_4_4_4_P(31),
  P(32) => R1IN_4_4_4_P(32),
  P(33) => R1IN_4_4_4_P(33),
  P(34) => R1IN_4_4_4_P(34),
  P(35) => R1IN_4_4_4_P(35),
  P(36) => R1IN_4_4_4_P(36),
  P(37) => R1IN_4_4_4_P(37),
  P(38) => R1IN_4_4_4_P(38),
  P(39) => R1IN_4_4_4_P(39),
  P(40) => R1IN_4_4_4_P(40),
  P(41) => R1IN_4_4_4_P(41),
  P(42) => R1IN_4_4_4_P(42),
  P(43) => R1IN_4_4_4_P(43),
  P(44) => R1IN_4_4_4_P(44),
  P(45) => R1IN_4_4_4_P(45),
  P(46) => R1IN_4_4_4_P(46),
  P(47) => R1IN_4_4_4_P(47),
  PCOUT(0) => R1IN_4_4_4_PCOUT(0),
  PCOUT(1) => R1IN_4_4_4_PCOUT(1),
  PCOUT(2) => R1IN_4_4_4_PCOUT(2),
  PCOUT(3) => R1IN_4_4_4_PCOUT(3),
  PCOUT(4) => R1IN_4_4_4_PCOUT(4),
  PCOUT(5) => R1IN_4_4_4_PCOUT(5),
  PCOUT(6) => R1IN_4_4_4_PCOUT(6),
  PCOUT(7) => R1IN_4_4_4_PCOUT(7),
  PCOUT(8) => R1IN_4_4_4_PCOUT(8),
  PCOUT(9) => R1IN_4_4_4_PCOUT(9),
  PCOUT(10) => R1IN_4_4_4_PCOUT(10),
  PCOUT(11) => R1IN_4_4_4_PCOUT(11),
  PCOUT(12) => R1IN_4_4_4_PCOUT(12),
  PCOUT(13) => R1IN_4_4_4_PCOUT(13),
  PCOUT(14) => R1IN_4_4_4_PCOUT(14),
  PCOUT(15) => R1IN_4_4_4_PCOUT(15),
  PCOUT(16) => R1IN_4_4_4_PCOUT(16),
  PCOUT(17) => R1IN_4_4_4_PCOUT(17),
  PCOUT(18) => R1IN_4_4_4_PCOUT(18),
  PCOUT(19) => R1IN_4_4_4_PCOUT(19),
  PCOUT(20) => R1IN_4_4_4_PCOUT(20),
  PCOUT(21) => R1IN_4_4_4_PCOUT(21),
  PCOUT(22) => R1IN_4_4_4_PCOUT(22),
  PCOUT(23) => R1IN_4_4_4_PCOUT(23),
  PCOUT(24) => R1IN_4_4_4_PCOUT(24),
  PCOUT(25) => R1IN_4_4_4_PCOUT(25),
  PCOUT(26) => R1IN_4_4_4_PCOUT(26),
  PCOUT(27) => R1IN_4_4_4_PCOUT(27),
  PCOUT(28) => R1IN_4_4_4_PCOUT(28),
  PCOUT(29) => R1IN_4_4_4_PCOUT(29),
  PCOUT(30) => R1IN_4_4_4_PCOUT(30),
  PCOUT(31) => R1IN_4_4_4_PCOUT(31),
  PCOUT(32) => R1IN_4_4_4_PCOUT(32),
  PCOUT(33) => R1IN_4_4_4_PCOUT(33),
  PCOUT(34) => R1IN_4_4_4_PCOUT(34),
  PCOUT(35) => R1IN_4_4_4_PCOUT(35),
  PCOUT(36) => R1IN_4_4_4_PCOUT(36),
  PCOUT(37) => R1IN_4_4_4_PCOUT(37),
  PCOUT(38) => R1IN_4_4_4_PCOUT(38),
  PCOUT(39) => R1IN_4_4_4_PCOUT(39),
  PCOUT(40) => R1IN_4_4_4_PCOUT(40),
  PCOUT(41) => R1IN_4_4_4_PCOUT(41),
  PCOUT(42) => R1IN_4_4_4_PCOUT(42),
  PCOUT(43) => R1IN_4_4_4_PCOUT(43),
  PCOUT(44) => R1IN_4_4_4_PCOUT(44),
  PCOUT(45) => R1IN_4_4_4_PCOUT(45),
  PCOUT(46) => R1IN_4_4_4_PCOUT(46),
  PCOUT(47) => R1IN_4_4_4_PCOUT(47));
R1IN_4_4_1q330w: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 0,
  MREG => 1,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18S"
)
port map (
  A(0) => A(34),
  A(1) => A(35),
  A(2) => A(36),
  A(3) => A(37),
  A(4) => A(38),
  A(5) => A(39),
  A(6) => A(40),
  A(7) => A(41),
  A(8) => A(42),
  A(9) => A(43),
  A(10) => A(44),
  A(11) => A(45),
  A(12) => A(46),
  A(13) => A(47),
  A(14) => A(48),
  A(15) => A(49),
  A(16) => A(50),
  A(17) => NN_1,
  B(0) => B(34),
  B(1) => B(35),
  B(2) => B(36),
  B(3) => B(37),
  B(4) => B(38),
  B(5) => B(39),
  B(6) => B(40),
  B(7) => B(41),
  B(8) => B(42),
  B(9) => B(43),
  B(10) => B(44),
  B(11) => B(45),
  B(12) => B(46),
  B(13) => B(47),
  B(14) => B(48),
  B(15) => B(49),
  B(16) => B(50),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => NN_1,
  PCIN(1) => NN_1,
  PCIN(2) => NN_1,
  PCIN(3) => NN_1,
  PCIN(4) => NN_1,
  PCIN(5) => NN_1,
  PCIN(6) => NN_1,
  PCIN(7) => NN_1,
  PCIN(8) => NN_1,
  PCIN(9) => NN_1,
  PCIN(10) => NN_1,
  PCIN(11) => NN_1,
  PCIN(12) => NN_1,
  PCIN(13) => NN_1,
  PCIN(14) => NN_1,
  PCIN(15) => NN_1,
  PCIN(16) => NN_1,
  PCIN(17) => NN_1,
  PCIN(18) => NN_1,
  PCIN(19) => NN_1,
  PCIN(20) => NN_1,
  PCIN(21) => NN_1,
  PCIN(22) => NN_1,
  PCIN(23) => NN_1,
  PCIN(24) => NN_1,
  PCIN(25) => NN_1,
  PCIN(26) => NN_1,
  PCIN(27) => NN_1,
  PCIN(28) => NN_1,
  PCIN(29) => NN_1,
  PCIN(30) => NN_1,
  PCIN(31) => NN_1,
  PCIN(32) => NN_1,
  PCIN(33) => NN_1,
  PCIN(34) => NN_1,
  PCIN(35) => NN_1,
  PCIN(36) => NN_1,
  PCIN(37) => NN_1,
  PCIN(38) => NN_1,
  PCIN(39) => NN_1,
  PCIN(40) => NN_1,
  PCIN(41) => NN_1,
  PCIN(42) => NN_1,
  PCIN(43) => NN_1,
  PCIN(44) => NN_1,
  PCIN(45) => NN_1,
  PCIN(46) => NN_1,
  PCIN(47) => NN_1,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_1,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => CLK,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => NN_1,
  CEM => EN,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_4_4_1_BCOUT(0),
  BCOUT(1) => R1IN_4_4_1_BCOUT(1),
  BCOUT(2) => R1IN_4_4_1_BCOUT(2),
  BCOUT(3) => R1IN_4_4_1_BCOUT(3),
  BCOUT(4) => R1IN_4_4_1_BCOUT(4),
  BCOUT(5) => R1IN_4_4_1_BCOUT(5),
  BCOUT(6) => R1IN_4_4_1_BCOUT(6),
  BCOUT(7) => R1IN_4_4_1_BCOUT(7),
  BCOUT(8) => R1IN_4_4_1_BCOUT(8),
  BCOUT(9) => R1IN_4_4_1_BCOUT(9),
  BCOUT(10) => R1IN_4_4_1_BCOUT(10),
  BCOUT(11) => R1IN_4_4_1_BCOUT(11),
  BCOUT(12) => R1IN_4_4_1_BCOUT(12),
  BCOUT(13) => R1IN_4_4_1_BCOUT(13),
  BCOUT(14) => R1IN_4_4_1_BCOUT(14),
  BCOUT(15) => R1IN_4_4_1_BCOUT(15),
  BCOUT(16) => R1IN_4_4_1_BCOUT(16),
  BCOUT(17) => R1IN_4_4_1_BCOUT(17),
  P(0) => R1IN_4_4F(0),
  P(1) => R1IN_4_4F(1),
  P(2) => R1IN_4_4F(2),
  P(3) => R1IN_4_4F(3),
  P(4) => R1IN_4_4F(4),
  P(5) => R1IN_4_4F(5),
  P(6) => R1IN_4_4F(6),
  P(7) => R1IN_4_4F(7),
  P(8) => R1IN_4_4F(8),
  P(9) => R1IN_4_4F(9),
  P(10) => R1IN_4_4F(10),
  P(11) => R1IN_4_4F(11),
  P(12) => R1IN_4_4F(12),
  P(13) => R1IN_4_4F(13),
  P(14) => R1IN_4_4F(14),
  P(15) => R1IN_4_4F(15),
  P(16) => R1IN_4_4F(16),
  P(17) => R1IN_4_4_ADD_2,
  P(18) => R1IN_4_4_1F(18),
  P(19) => R1IN_4_4_1F(19),
  P(20) => R1IN_4_4_1F(20),
  P(21) => R1IN_4_4_1F(21),
  P(22) => R1IN_4_4_1F(22),
  P(23) => R1IN_4_4_1F(23),
  P(24) => R1IN_4_4_1F(24),
  P(25) => R1IN_4_4_1F(25),
  P(26) => R1IN_4_4_1F(26),
  P(27) => R1IN_4_4_1F(27),
  P(28) => R1IN_4_4_1F(28),
  P(29) => R1IN_4_4_1F(29),
  P(30) => R1IN_4_4_1F(30),
  P(31) => R1IN_4_4_1F(31),
  P(32) => R1IN_4_4_1F(32),
  P(33) => R1IN_4_4_1F(33),
  P(34) => UC_236,
  P(35) => UC_237,
  P(36) => UC_238,
  P(37) => UC_239,
  P(38) => UC_240,
  P(39) => UC_241,
  P(40) => UC_242,
  P(41) => UC_243,
  P(42) => UC_244,
  P(43) => UC_245,
  P(44) => UC_246,
  P(45) => UC_247,
  P(46) => UC_248,
  P(47) => UC_249,
  PCOUT(0) => R1IN_4_4_1_PCOUT(0),
  PCOUT(1) => R1IN_4_4_1_PCOUT(1),
  PCOUT(2) => R1IN_4_4_1_PCOUT(2),
  PCOUT(3) => R1IN_4_4_1_PCOUT(3),
  PCOUT(4) => R1IN_4_4_1_PCOUT(4),
  PCOUT(5) => R1IN_4_4_1_PCOUT(5),
  PCOUT(6) => R1IN_4_4_1_PCOUT(6),
  PCOUT(7) => R1IN_4_4_1_PCOUT(7),
  PCOUT(8) => R1IN_4_4_1_PCOUT(8),
  PCOUT(9) => R1IN_4_4_1_PCOUT(9),
  PCOUT(10) => R1IN_4_4_1_PCOUT(10),
  PCOUT(11) => R1IN_4_4_1_PCOUT(11),
  PCOUT(12) => R1IN_4_4_1_PCOUT(12),
  PCOUT(13) => R1IN_4_4_1_PCOUT(13),
  PCOUT(14) => R1IN_4_4_1_PCOUT(14),
  PCOUT(15) => R1IN_4_4_1_PCOUT(15),
  PCOUT(16) => R1IN_4_4_1_PCOUT(16),
  PCOUT(17) => R1IN_4_4_1_PCOUT(17),
  PCOUT(18) => R1IN_4_4_1_PCOUT(18),
  PCOUT(19) => R1IN_4_4_1_PCOUT(19),
  PCOUT(20) => R1IN_4_4_1_PCOUT(20),
  PCOUT(21) => R1IN_4_4_1_PCOUT(21),
  PCOUT(22) => R1IN_4_4_1_PCOUT(22),
  PCOUT(23) => R1IN_4_4_1_PCOUT(23),
  PCOUT(24) => R1IN_4_4_1_PCOUT(24),
  PCOUT(25) => R1IN_4_4_1_PCOUT(25),
  PCOUT(26) => R1IN_4_4_1_PCOUT(26),
  PCOUT(27) => R1IN_4_4_1_PCOUT(27),
  PCOUT(28) => R1IN_4_4_1_PCOUT(28),
  PCOUT(29) => R1IN_4_4_1_PCOUT(29),
  PCOUT(30) => R1IN_4_4_1_PCOUT(30),
  PCOUT(31) => R1IN_4_4_1_PCOUT(31),
  PCOUT(32) => R1IN_4_4_1_PCOUT(32),
  PCOUT(33) => R1IN_4_4_1_PCOUT(33),
  PCOUT(34) => R1IN_4_4_1_PCOUT(34),
  PCOUT(35) => R1IN_4_4_1_PCOUT(35),
  PCOUT(36) => R1IN_4_4_1_PCOUT(36),
  PCOUT(37) => R1IN_4_4_1_PCOUT(37),
  PCOUT(38) => R1IN_4_4_1_PCOUT(38),
  PCOUT(39) => R1IN_4_4_1_PCOUT(39),
  PCOUT(40) => R1IN_4_4_1_PCOUT(40),
  PCOUT(41) => R1IN_4_4_1_PCOUT(41),
  PCOUT(42) => R1IN_4_4_1_PCOUT(42),
  PCOUT(43) => R1IN_4_4_1_PCOUT(43),
  PCOUT(44) => R1IN_4_4_1_PCOUT(44),
  PCOUT(45) => R1IN_4_4_1_PCOUT(45),
  PCOUT(46) => R1IN_4_4_1_PCOUT(46),
  PCOUT(47) => R1IN_4_4_1_PCOUT(47));
R1IN_4_1q330w: DSP48 
generic map(
  AREG => 1,
  BREG => 1,
  CREG => 0,
  PREG => 1,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => A(17),
  A(1) => A(18),
  A(2) => A(19),
  A(3) => A(20),
  A(4) => A(21),
  A(5) => A(22),
  A(6) => A(23),
  A(7) => A(24),
  A(8) => A(25),
  A(9) => A(26),
  A(10) => A(27),
  A(11) => A(28),
  A(12) => A(29),
  A(13) => A(30),
  A(14) => A(31),
  A(15) => A(32),
  A(16) => A(33),
  A(17) => NN_1,
  B(0) => B(17),
  B(1) => B(18),
  B(2) => B(19),
  B(3) => B(20),
  B(4) => B(21),
  B(5) => B(22),
  B(6) => B(23),
  B(7) => B(24),
  B(8) => B(25),
  B(9) => B(26),
  B(10) => B(27),
  B(11) => B(28),
  B(12) => B(29),
  B(13) => B(30),
  B(14) => B(31),
  B(15) => B(32),
  B(16) => B(33),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => NN_1,
  PCIN(1) => NN_1,
  PCIN(2) => NN_1,
  PCIN(3) => NN_1,
  PCIN(4) => NN_1,
  PCIN(5) => NN_1,
  PCIN(6) => NN_1,
  PCIN(7) => NN_1,
  PCIN(8) => NN_1,
  PCIN(9) => NN_1,
  PCIN(10) => NN_1,
  PCIN(11) => NN_1,
  PCIN(12) => NN_1,
  PCIN(13) => NN_1,
  PCIN(14) => NN_1,
  PCIN(15) => NN_1,
  PCIN(16) => NN_1,
  PCIN(17) => NN_1,
  PCIN(18) => NN_1,
  PCIN(19) => NN_1,
  PCIN(20) => NN_1,
  PCIN(21) => NN_1,
  PCIN(22) => NN_1,
  PCIN(23) => NN_1,
  PCIN(24) => NN_1,
  PCIN(25) => NN_1,
  PCIN(26) => NN_1,
  PCIN(27) => NN_1,
  PCIN(28) => NN_1,
  PCIN(29) => NN_1,
  PCIN(30) => NN_1,
  PCIN(31) => NN_1,
  PCIN(32) => NN_1,
  PCIN(33) => NN_1,
  PCIN(34) => NN_1,
  PCIN(35) => NN_1,
  PCIN(36) => NN_1,
  PCIN(37) => NN_1,
  PCIN(38) => NN_1,
  PCIN(39) => NN_1,
  PCIN(40) => NN_1,
  PCIN(41) => NN_1,
  PCIN(42) => NN_1,
  PCIN(43) => NN_1,
  PCIN(44) => NN_1,
  PCIN(45) => NN_1,
  PCIN(46) => NN_1,
  PCIN(47) => NN_1,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_1,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => CLK,
  CEA => EN,
  CEB => EN,
  CEC => NN_1,
  CEP => EN,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_4_1_BCOUT(0),
  BCOUT(1) => R1IN_4_1_BCOUT(1),
  BCOUT(2) => R1IN_4_1_BCOUT(2),
  BCOUT(3) => R1IN_4_1_BCOUT(3),
  BCOUT(4) => R1IN_4_1_BCOUT(4),
  BCOUT(5) => R1IN_4_1_BCOUT(5),
  BCOUT(6) => R1IN_4_1_BCOUT(6),
  BCOUT(7) => R1IN_4_1_BCOUT(7),
  BCOUT(8) => R1IN_4_1_BCOUT(8),
  BCOUT(9) => R1IN_4_1_BCOUT(9),
  BCOUT(10) => R1IN_4_1_BCOUT(10),
  BCOUT(11) => R1IN_4_1_BCOUT(11),
  BCOUT(12) => R1IN_4_1_BCOUT(12),
  BCOUT(13) => R1IN_4_1_BCOUT(13),
  BCOUT(14) => R1IN_4_1_BCOUT(14),
  BCOUT(15) => R1IN_4_1_BCOUT(15),
  BCOUT(16) => R1IN_4_1_BCOUT(16),
  BCOUT(17) => R1IN_4_1_BCOUT(17),
  P(0) => R1IN_4FF(0),
  P(1) => R1IN_4FF(1),
  P(2) => R1IN_4FF(2),
  P(3) => R1IN_4FF(3),
  P(4) => R1IN_4FF(4),
  P(5) => R1IN_4FF(5),
  P(6) => R1IN_4FF(6),
  P(7) => R1IN_4FF(7),
  P(8) => R1IN_4FF(8),
  P(9) => R1IN_4FF(9),
  P(10) => R1IN_4FF(10),
  P(11) => R1IN_4FF(11),
  P(12) => R1IN_4FF(12),
  P(13) => R1IN_4FF(13),
  P(14) => R1IN_4FF(14),
  P(15) => R1IN_4FF(15),
  P(16) => R1IN_4FF(16),
  P(17) => R1IN_4_1F_RETO(17),
  P(18) => R1IN_4_1F_RETO(18),
  P(19) => R1IN_4_1F_RETO(19),
  P(20) => R1IN_4_1F_RETO(20),
  P(21) => R1IN_4_1F_RETO(21),
  P(22) => R1IN_4_1F_RETO(22),
  P(23) => R1IN_4_1F_RETO(23),
  P(24) => R1IN_4_1F_RETO(24),
  P(25) => R1IN_4_1F_RETO(25),
  P(26) => R1IN_4_1F_RETO(26),
  P(27) => R1IN_4_1F_RETO(27),
  P(28) => R1IN_4_1F_RETO(28),
  P(29) => R1IN_4_1F_RETO(29),
  P(30) => R1IN_4_1F_RETO(30),
  P(31) => R1IN_4_1F_RETO(31),
  P(32) => R1IN_4_1F_RETO(32),
  P(33) => R1IN_4_1F_RETO(33),
  P(34) => R1IN_4_1_P(34),
  P(35) => R1IN_4_1_P(35),
  P(36) => R1IN_4_1_P(36),
  P(37) => R1IN_4_1_P(37),
  P(38) => R1IN_4_1_P(38),
  P(39) => R1IN_4_1_P(39),
  P(40) => R1IN_4_1_P(40),
  P(41) => R1IN_4_1_P(41),
  P(42) => R1IN_4_1_P(42),
  P(43) => R1IN_4_1_P(43),
  P(44) => R1IN_4_1_P(44),
  P(45) => R1IN_4_1_P(45),
  P(46) => R1IN_4_1_P(46),
  P(47) => R1IN_4_1_P(47),
  PCOUT(0) => R1IN_4_1_PCOUT(0),
  PCOUT(1) => R1IN_4_1_PCOUT(1),
  PCOUT(2) => R1IN_4_1_PCOUT(2),
  PCOUT(3) => R1IN_4_1_PCOUT(3),
  PCOUT(4) => R1IN_4_1_PCOUT(4),
  PCOUT(5) => R1IN_4_1_PCOUT(5),
  PCOUT(6) => R1IN_4_1_PCOUT(6),
  PCOUT(7) => R1IN_4_1_PCOUT(7),
  PCOUT(8) => R1IN_4_1_PCOUT(8),
  PCOUT(9) => R1IN_4_1_PCOUT(9),
  PCOUT(10) => R1IN_4_1_PCOUT(10),
  PCOUT(11) => R1IN_4_1_PCOUT(11),
  PCOUT(12) => R1IN_4_1_PCOUT(12),
  PCOUT(13) => R1IN_4_1_PCOUT(13),
  PCOUT(14) => R1IN_4_1_PCOUT(14),
  PCOUT(15) => R1IN_4_1_PCOUT(15),
  PCOUT(16) => R1IN_4_1_PCOUT(16),
  PCOUT(17) => R1IN_4_1_PCOUT(17),
  PCOUT(18) => R1IN_4_1_PCOUT(18),
  PCOUT(19) => R1IN_4_1_PCOUT(19),
  PCOUT(20) => R1IN_4_1_PCOUT(20),
  PCOUT(21) => R1IN_4_1_PCOUT(21),
  PCOUT(22) => R1IN_4_1_PCOUT(22),
  PCOUT(23) => R1IN_4_1_PCOUT(23),
  PCOUT(24) => R1IN_4_1_PCOUT(24),
  PCOUT(25) => R1IN_4_1_PCOUT(25),
  PCOUT(26) => R1IN_4_1_PCOUT(26),
  PCOUT(27) => R1IN_4_1_PCOUT(27),
  PCOUT(28) => R1IN_4_1_PCOUT(28),
  PCOUT(29) => R1IN_4_1_PCOUT(29),
  PCOUT(30) => R1IN_4_1_PCOUT(30),
  PCOUT(31) => R1IN_4_1_PCOUT(31),
  PCOUT(32) => R1IN_4_1_PCOUT(32),
  PCOUT(33) => R1IN_4_1_PCOUT(33),
  PCOUT(34) => R1IN_4_1_PCOUT(34),
  PCOUT(35) => R1IN_4_1_PCOUT(35),
  PCOUT(36) => R1IN_4_1_PCOUT(36),
  PCOUT(37) => R1IN_4_1_PCOUT(37),
  PCOUT(38) => R1IN_4_1_PCOUT(38),
  PCOUT(39) => R1IN_4_1_PCOUT(39),
  PCOUT(40) => R1IN_4_1_PCOUT(40),
  PCOUT(41) => R1IN_4_1_PCOUT(41),
  PCOUT(42) => R1IN_4_1_PCOUT(42),
  PCOUT(43) => R1IN_4_1_PCOUT(43),
  PCOUT(44) => R1IN_4_1_PCOUT(44),
  PCOUT(45) => R1IN_4_1_PCOUT(45),
  PCOUT(46) => R1IN_4_1_PCOUT(46),
  PCOUT(47) => R1IN_4_1_PCOUT(47));
R1IN_3_1q330w: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 0,
  MREG => 1,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18S"
)
port map (
  A(0) => B(17),
  A(1) => B(18),
  A(2) => B(19),
  A(3) => B(20),
  A(4) => B(21),
  A(5) => B(22),
  A(6) => B(23),
  A(7) => B(24),
  A(8) => B(25),
  A(9) => B(26),
  A(10) => B(27),
  A(11) => B(28),
  A(12) => B(29),
  A(13) => B(30),
  A(14) => B(31),
  A(15) => B(32),
  A(16) => B(33),
  A(17) => NN_1,
  B(0) => A(0),
  B(1) => A(1),
  B(2) => A(2),
  B(3) => A(3),
  B(4) => A(4),
  B(5) => A(5),
  B(6) => A(6),
  B(7) => A(7),
  B(8) => A(8),
  B(9) => A(9),
  B(10) => A(10),
  B(11) => A(11),
  B(12) => A(12),
  B(13) => A(13),
  B(14) => A(14),
  B(15) => A(15),
  B(16) => A(16),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => NN_1,
  PCIN(1) => NN_1,
  PCIN(2) => NN_1,
  PCIN(3) => NN_1,
  PCIN(4) => NN_1,
  PCIN(5) => NN_1,
  PCIN(6) => NN_1,
  PCIN(7) => NN_1,
  PCIN(8) => NN_1,
  PCIN(9) => NN_1,
  PCIN(10) => NN_1,
  PCIN(11) => NN_1,
  PCIN(12) => NN_1,
  PCIN(13) => NN_1,
  PCIN(14) => NN_1,
  PCIN(15) => NN_1,
  PCIN(16) => NN_1,
  PCIN(17) => NN_1,
  PCIN(18) => NN_1,
  PCIN(19) => NN_1,
  PCIN(20) => NN_1,
  PCIN(21) => NN_1,
  PCIN(22) => NN_1,
  PCIN(23) => NN_1,
  PCIN(24) => NN_1,
  PCIN(25) => NN_1,
  PCIN(26) => NN_1,
  PCIN(27) => NN_1,
  PCIN(28) => NN_1,
  PCIN(29) => NN_1,
  PCIN(30) => NN_1,
  PCIN(31) => NN_1,
  PCIN(32) => NN_1,
  PCIN(33) => NN_1,
  PCIN(34) => NN_1,
  PCIN(35) => NN_1,
  PCIN(36) => NN_1,
  PCIN(37) => NN_1,
  PCIN(38) => NN_1,
  PCIN(39) => NN_1,
  PCIN(40) => NN_1,
  PCIN(41) => NN_1,
  PCIN(42) => NN_1,
  PCIN(43) => NN_1,
  PCIN(44) => NN_1,
  PCIN(45) => NN_1,
  PCIN(46) => NN_1,
  PCIN(47) => NN_1,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_1,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => CLK,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => NN_1,
  CEM => EN,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_3_1_BCOUT(0),
  BCOUT(1) => R1IN_3_1_BCOUT(1),
  BCOUT(2) => R1IN_3_1_BCOUT(2),
  BCOUT(3) => R1IN_3_1_BCOUT(3),
  BCOUT(4) => R1IN_3_1_BCOUT(4),
  BCOUT(5) => R1IN_3_1_BCOUT(5),
  BCOUT(6) => R1IN_3_1_BCOUT(6),
  BCOUT(7) => R1IN_3_1_BCOUT(7),
  BCOUT(8) => R1IN_3_1_BCOUT(8),
  BCOUT(9) => R1IN_3_1_BCOUT(9),
  BCOUT(10) => R1IN_3_1_BCOUT(10),
  BCOUT(11) => R1IN_3_1_BCOUT(11),
  BCOUT(12) => R1IN_3_1_BCOUT(12),
  BCOUT(13) => R1IN_3_1_BCOUT(13),
  BCOUT(14) => R1IN_3_1_BCOUT(14),
  BCOUT(15) => R1IN_3_1_BCOUT(15),
  BCOUT(16) => R1IN_3_1_BCOUT(16),
  BCOUT(17) => R1IN_3_1_BCOUT(17),
  P(0) => R1IN_3F(0),
  P(1) => R1IN_3F(1),
  P(2) => R1IN_3F(2),
  P(3) => R1IN_3F(3),
  P(4) => R1IN_3F(4),
  P(5) => R1IN_3F(5),
  P(6) => R1IN_3F(6),
  P(7) => R1IN_3F(7),
  P(8) => R1IN_3F(8),
  P(9) => R1IN_3F(9),
  P(10) => R1IN_3F(10),
  P(11) => R1IN_3F(11),
  P(12) => R1IN_3F(12),
  P(13) => R1IN_3F(13),
  P(14) => R1IN_3F(14),
  P(15) => R1IN_3F(15),
  P(16) => R1IN_3F(16),
  P(17) => R1IN_3_1F(17),
  P(18) => R1IN_3_1F(18),
  P(19) => R1IN_3_1F(19),
  P(20) => R1IN_3_1F(20),
  P(21) => R1IN_3_1F(21),
  P(22) => R1IN_3_1F(22),
  P(23) => R1IN_3_1F(23),
  P(24) => R1IN_3_1F(24),
  P(25) => R1IN_3_1F(25),
  P(26) => R1IN_3_1F(26),
  P(27) => R1IN_3_1F(27),
  P(28) => R1IN_3_1F(28),
  P(29) => R1IN_3_1F(29),
  P(30) => R1IN_3_1F(30),
  P(31) => R1IN_3_1F(31),
  P(32) => R1IN_3_1F(32),
  P(33) => R1IN_3_1F(33),
  P(34) => UC_208,
  P(35) => UC_209,
  P(36) => UC_210,
  P(37) => UC_211,
  P(38) => UC_212,
  P(39) => UC_213,
  P(40) => UC_214,
  P(41) => UC_215,
  P(42) => UC_216,
  P(43) => UC_217,
  P(44) => UC_218,
  P(45) => UC_219,
  P(46) => UC_220,
  P(47) => UC_221,
  PCOUT(0) => R1IN_3_1_PCOUT(0),
  PCOUT(1) => R1IN_3_1_PCOUT(1),
  PCOUT(2) => R1IN_3_1_PCOUT(2),
  PCOUT(3) => R1IN_3_1_PCOUT(3),
  PCOUT(4) => R1IN_3_1_PCOUT(4),
  PCOUT(5) => R1IN_3_1_PCOUT(5),
  PCOUT(6) => R1IN_3_1_PCOUT(6),
  PCOUT(7) => R1IN_3_1_PCOUT(7),
  PCOUT(8) => R1IN_3_1_PCOUT(8),
  PCOUT(9) => R1IN_3_1_PCOUT(9),
  PCOUT(10) => R1IN_3_1_PCOUT(10),
  PCOUT(11) => R1IN_3_1_PCOUT(11),
  PCOUT(12) => R1IN_3_1_PCOUT(12),
  PCOUT(13) => R1IN_3_1_PCOUT(13),
  PCOUT(14) => R1IN_3_1_PCOUT(14),
  PCOUT(15) => R1IN_3_1_PCOUT(15),
  PCOUT(16) => R1IN_3_1_PCOUT(16),
  PCOUT(17) => R1IN_3_1_PCOUT(17),
  PCOUT(18) => R1IN_3_1_PCOUT(18),
  PCOUT(19) => R1IN_3_1_PCOUT(19),
  PCOUT(20) => R1IN_3_1_PCOUT(20),
  PCOUT(21) => R1IN_3_1_PCOUT(21),
  PCOUT(22) => R1IN_3_1_PCOUT(22),
  PCOUT(23) => R1IN_3_1_PCOUT(23),
  PCOUT(24) => R1IN_3_1_PCOUT(24),
  PCOUT(25) => R1IN_3_1_PCOUT(25),
  PCOUT(26) => R1IN_3_1_PCOUT(26),
  PCOUT(27) => R1IN_3_1_PCOUT(27),
  PCOUT(28) => R1IN_3_1_PCOUT(28),
  PCOUT(29) => R1IN_3_1_PCOUT(29),
  PCOUT(30) => R1IN_3_1_PCOUT(30),
  PCOUT(31) => R1IN_3_1_PCOUT(31),
  PCOUT(32) => R1IN_3_1_PCOUT(32),
  PCOUT(33) => R1IN_3_1_PCOUT(33),
  PCOUT(34) => R1IN_3_1_PCOUT(34),
  PCOUT(35) => R1IN_3_1_PCOUT(35),
  PCOUT(36) => R1IN_3_1_PCOUT(36),
  PCOUT(37) => R1IN_3_1_PCOUT(37),
  PCOUT(38) => R1IN_3_1_PCOUT(38),
  PCOUT(39) => R1IN_3_1_PCOUT(39),
  PCOUT(40) => R1IN_3_1_PCOUT(40),
  PCOUT(41) => R1IN_3_1_PCOUT(41),
  PCOUT(42) => R1IN_3_1_PCOUT(42),
  PCOUT(43) => R1IN_3_1_PCOUT(43),
  PCOUT(44) => R1IN_3_1_PCOUT(44),
  PCOUT(45) => R1IN_3_1_PCOUT(45),
  PCOUT(46) => R1IN_3_1_PCOUT(46),
  PCOUT(47) => R1IN_3_1_PCOUT(47));
R1IN_2_1q330w: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 1,
  MREG => 1,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18S"
)
port map (
  A(0) => A(17),
  A(1) => A(18),
  A(2) => A(19),
  A(3) => A(20),
  A(4) => A(21),
  A(5) => A(22),
  A(6) => A(23),
  A(7) => A(24),
  A(8) => A(25),
  A(9) => A(26),
  A(10) => A(27),
  A(11) => A(28),
  A(12) => A(29),
  A(13) => A(30),
  A(14) => A(31),
  A(15) => A(32),
  A(16) => A(33),
  A(17) => NN_1,
  B(0) => B(0),
  B(1) => B(1),
  B(2) => B(2),
  B(3) => B(3),
  B(4) => B(4),
  B(5) => B(5),
  B(6) => B(6),
  B(7) => B(7),
  B(8) => B(8),
  B(9) => B(9),
  B(10) => B(10),
  B(11) => B(11),
  B(12) => B(12),
  B(13) => B(13),
  B(14) => B(14),
  B(15) => B(15),
  B(16) => B(16),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => NN_1,
  PCIN(1) => NN_1,
  PCIN(2) => NN_1,
  PCIN(3) => NN_1,
  PCIN(4) => NN_1,
  PCIN(5) => NN_1,
  PCIN(6) => NN_1,
  PCIN(7) => NN_1,
  PCIN(8) => NN_1,
  PCIN(9) => NN_1,
  PCIN(10) => NN_1,
  PCIN(11) => NN_1,
  PCIN(12) => NN_1,
  PCIN(13) => NN_1,
  PCIN(14) => NN_1,
  PCIN(15) => NN_1,
  PCIN(16) => NN_1,
  PCIN(17) => NN_1,
  PCIN(18) => NN_1,
  PCIN(19) => NN_1,
  PCIN(20) => NN_1,
  PCIN(21) => NN_1,
  PCIN(22) => NN_1,
  PCIN(23) => NN_1,
  PCIN(24) => NN_1,
  PCIN(25) => NN_1,
  PCIN(26) => NN_1,
  PCIN(27) => NN_1,
  PCIN(28) => NN_1,
  PCIN(29) => NN_1,
  PCIN(30) => NN_1,
  PCIN(31) => NN_1,
  PCIN(32) => NN_1,
  PCIN(33) => NN_1,
  PCIN(34) => NN_1,
  PCIN(35) => NN_1,
  PCIN(36) => NN_1,
  PCIN(37) => NN_1,
  PCIN(38) => NN_1,
  PCIN(39) => NN_1,
  PCIN(40) => NN_1,
  PCIN(41) => NN_1,
  PCIN(42) => NN_1,
  PCIN(43) => NN_1,
  PCIN(44) => NN_1,
  PCIN(45) => NN_1,
  PCIN(46) => NN_1,
  PCIN(47) => NN_1,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_1,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => CLK,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => EN,
  CEM => EN,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => B_0(0),
  BCOUT(1) => B_0(1),
  BCOUT(2) => B_0(2),
  BCOUT(3) => B_0(3),
  BCOUT(4) => B_0(4),
  BCOUT(5) => B_0(5),
  BCOUT(6) => B_0(6),
  BCOUT(7) => B_0(7),
  BCOUT(8) => B_0(8),
  BCOUT(9) => B_0(9),
  BCOUT(10) => B_0(10),
  BCOUT(11) => B_0(11),
  BCOUT(12) => B_0(12),
  BCOUT(13) => B_0(13),
  BCOUT(14) => B_0(14),
  BCOUT(15) => B_0(15),
  BCOUT(16) => B_0(16),
  BCOUT(17) => GND_0,
  P(0) => R1IN_2F_RETO(0),
  P(1) => R1IN_2F_RETO(1),
  P(2) => R1IN_2F_RETO(2),
  P(3) => R1IN_2F_RETO(3),
  P(4) => R1IN_2F_RETO(4),
  P(5) => R1IN_2F_RETO(5),
  P(6) => R1IN_2F_RETO(6),
  P(7) => R1IN_2F_RETO(7),
  P(8) => R1IN_2F_RETO(8),
  P(9) => R1IN_2F_RETO(9),
  P(10) => R1IN_2F_RETO(10),
  P(11) => R1IN_2F_RETO(11),
  P(12) => R1IN_2F_RETO(12),
  P(13) => R1IN_2F_RETO(13),
  P(14) => R1IN_2F_RETO(14),
  P(15) => R1IN_2F_RETO(15),
  P(16) => R1IN_2F_RETO(16),
  P(17) => R1IN_2_1F_RETO(17),
  P(18) => R1IN_2_1F_RETO(18),
  P(19) => R1IN_2_1F_RETO(19),
  P(20) => R1IN_2_1F_RETO(20),
  P(21) => R1IN_2_1F_RETO(21),
  P(22) => R1IN_2_1F_RETO(22),
  P(23) => R1IN_2_1F_RETO(23),
  P(24) => R1IN_2_1F_RETO(24),
  P(25) => R1IN_2_1F_RETO(25),
  P(26) => R1IN_2_1F_RETO(26),
  P(27) => R1IN_2_1F_RETO(27),
  P(28) => R1IN_2_1F_RETO(28),
  P(29) => R1IN_2_1F_RETO(29),
  P(30) => R1IN_2_1F_RETO(30),
  P(31) => R1IN_2_1F_RETO(31),
  P(32) => R1IN_2_1F_RETO(32),
  P(33) => R1IN_2_1F_RETO(33),
  P(34) => R1IN_2_1_P(34),
  P(35) => R1IN_2_1_P(35),
  P(36) => R1IN_2_1_P(36),
  P(37) => R1IN_2_1_P(37),
  P(38) => R1IN_2_1_P(38),
  P(39) => R1IN_2_1_P(39),
  P(40) => R1IN_2_1_P(40),
  P(41) => R1IN_2_1_P(41),
  P(42) => R1IN_2_1_P(42),
  P(43) => R1IN_2_1_P(43),
  P(44) => R1IN_2_1_P(44),
  P(45) => R1IN_2_1_P(45),
  P(46) => R1IN_2_1_P(46),
  P(47) => R1IN_2_1_P(47),
  PCOUT(0) => R1IN_2_1_PCOUT(0),
  PCOUT(1) => R1IN_2_1_PCOUT(1),
  PCOUT(2) => R1IN_2_1_PCOUT(2),
  PCOUT(3) => R1IN_2_1_PCOUT(3),
  PCOUT(4) => R1IN_2_1_PCOUT(4),
  PCOUT(5) => R1IN_2_1_PCOUT(5),
  PCOUT(6) => R1IN_2_1_PCOUT(6),
  PCOUT(7) => R1IN_2_1_PCOUT(7),
  PCOUT(8) => R1IN_2_1_PCOUT(8),
  PCOUT(9) => R1IN_2_1_PCOUT(9),
  PCOUT(10) => R1IN_2_1_PCOUT(10),
  PCOUT(11) => R1IN_2_1_PCOUT(11),
  PCOUT(12) => R1IN_2_1_PCOUT(12),
  PCOUT(13) => R1IN_2_1_PCOUT(13),
  PCOUT(14) => R1IN_2_1_PCOUT(14),
  PCOUT(15) => R1IN_2_1_PCOUT(15),
  PCOUT(16) => R1IN_2_1_PCOUT(16),
  PCOUT(17) => R1IN_2_1_PCOUT(17),
  PCOUT(18) => R1IN_2_1_PCOUT(18),
  PCOUT(19) => R1IN_2_1_PCOUT(19),
  PCOUT(20) => R1IN_2_1_PCOUT(20),
  PCOUT(21) => R1IN_2_1_PCOUT(21),
  PCOUT(22) => R1IN_2_1_PCOUT(22),
  PCOUT(23) => R1IN_2_1_PCOUT(23),
  PCOUT(24) => R1IN_2_1_PCOUT(24),
  PCOUT(25) => R1IN_2_1_PCOUT(25),
  PCOUT(26) => R1IN_2_1_PCOUT(26),
  PCOUT(27) => R1IN_2_1_PCOUT(27),
  PCOUT(28) => R1IN_2_1_PCOUT(28),
  PCOUT(29) => R1IN_2_1_PCOUT(29),
  PCOUT(30) => R1IN_2_1_PCOUT(30),
  PCOUT(31) => R1IN_2_1_PCOUT(31),
  PCOUT(32) => R1IN_2_1_PCOUT(32),
  PCOUT(33) => R1IN_2_1_PCOUT(33),
  PCOUT(34) => R1IN_2_1_PCOUT(34),
  PCOUT(35) => R1IN_2_1_PCOUT(35),
  PCOUT(36) => R1IN_2_1_PCOUT(36),
  PCOUT(37) => R1IN_2_1_PCOUT(37),
  PCOUT(38) => R1IN_2_1_PCOUT(38),
  PCOUT(39) => R1IN_2_1_PCOUT(39),
  PCOUT(40) => R1IN_2_1_PCOUT(40),
  PCOUT(41) => R1IN_2_1_PCOUT(41),
  PCOUT(42) => R1IN_2_1_PCOUT(42),
  PCOUT(43) => R1IN_2_1_PCOUT(43),
  PCOUT(44) => R1IN_2_1_PCOUT(44),
  PCOUT(45) => R1IN_2_1_PCOUT(45),
  PCOUT(46) => R1IN_2_1_PCOUT(46),
  PCOUT(47) => R1IN_2_1_PCOUT(47));
R1IN_1q330w: DSP48 
generic map(
  AREG => 1,
  BREG => 1,
  CREG => 0,
  PREG => 1,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "CASCADE",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => A(0),
  A(1) => A(1),
  A(2) => A(2),
  A(3) => A(3),
  A(4) => A(4),
  A(5) => A(5),
  A(6) => A(6),
  A(7) => A(7),
  A(8) => A(8),
  A(9) => A(9),
  A(10) => A(10),
  A(11) => A(11),
  A(12) => A(12),
  A(13) => A(13),
  A(14) => A(14),
  A(15) => A(15),
  A(16) => A(16),
  A(17) => NN_1,
  B(0) => NN_1,
  B(1) => NN_1,
  B(2) => NN_1,
  B(3) => NN_1,
  B(4) => NN_1,
  B(5) => NN_1,
  B(6) => NN_1,
  B(7) => NN_1,
  B(8) => NN_1,
  B(9) => NN_1,
  B(10) => NN_1,
  B(11) => NN_1,
  B(12) => NN_1,
  B(13) => NN_1,
  B(14) => NN_1,
  B(15) => NN_1,
  B(16) => NN_1,
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => B_0(0),
  BCIN(1) => B_0(1),
  BCIN(2) => B_0(2),
  BCIN(3) => B_0(3),
  BCIN(4) => B_0(4),
  BCIN(5) => B_0(5),
  BCIN(6) => B_0(6),
  BCIN(7) => B_0(7),
  BCIN(8) => B_0(8),
  BCIN(9) => B_0(9),
  BCIN(10) => B_0(10),
  BCIN(11) => B_0(11),
  BCIN(12) => B_0(12),
  BCIN(13) => B_0(13),
  BCIN(14) => B_0(14),
  BCIN(15) => B_0(15),
  BCIN(16) => B_0(16),
  BCIN(17) => GND_0,
  PCIN(0) => NN_1,
  PCIN(1) => NN_1,
  PCIN(2) => NN_1,
  PCIN(3) => NN_1,
  PCIN(4) => NN_1,
  PCIN(5) => NN_1,
  PCIN(6) => NN_1,
  PCIN(7) => NN_1,
  PCIN(8) => NN_1,
  PCIN(9) => NN_1,
  PCIN(10) => NN_1,
  PCIN(11) => NN_1,
  PCIN(12) => NN_1,
  PCIN(13) => NN_1,
  PCIN(14) => NN_1,
  PCIN(15) => NN_1,
  PCIN(16) => NN_1,
  PCIN(17) => NN_1,
  PCIN(18) => NN_1,
  PCIN(19) => NN_1,
  PCIN(20) => NN_1,
  PCIN(21) => NN_1,
  PCIN(22) => NN_1,
  PCIN(23) => NN_1,
  PCIN(24) => NN_1,
  PCIN(25) => NN_1,
  PCIN(26) => NN_1,
  PCIN(27) => NN_1,
  PCIN(28) => NN_1,
  PCIN(29) => NN_1,
  PCIN(30) => NN_1,
  PCIN(31) => NN_1,
  PCIN(32) => NN_1,
  PCIN(33) => NN_1,
  PCIN(34) => NN_1,
  PCIN(35) => NN_1,
  PCIN(36) => NN_1,
  PCIN(37) => NN_1,
  PCIN(38) => NN_1,
  PCIN(39) => NN_1,
  PCIN(40) => NN_1,
  PCIN(41) => NN_1,
  PCIN(42) => NN_1,
  PCIN(43) => NN_1,
  PCIN(44) => NN_1,
  PCIN(45) => NN_1,
  PCIN(46) => NN_1,
  PCIN(47) => NN_1,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_1,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => CLK,
  CEA => EN,
  CEB => EN,
  CEC => NN_1,
  CEP => EN,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_1_BCOUT(0),
  BCOUT(1) => R1IN_1_BCOUT(1),
  BCOUT(2) => R1IN_1_BCOUT(2),
  BCOUT(3) => R1IN_1_BCOUT(3),
  BCOUT(4) => R1IN_1_BCOUT(4),
  BCOUT(5) => R1IN_1_BCOUT(5),
  BCOUT(6) => R1IN_1_BCOUT(6),
  BCOUT(7) => R1IN_1_BCOUT(7),
  BCOUT(8) => R1IN_1_BCOUT(8),
  BCOUT(9) => R1IN_1_BCOUT(9),
  BCOUT(10) => R1IN_1_BCOUT(10),
  BCOUT(11) => R1IN_1_BCOUT(11),
  BCOUT(12) => R1IN_1_BCOUT(12),
  BCOUT(13) => R1IN_1_BCOUT(13),
  BCOUT(14) => R1IN_1_BCOUT(14),
  BCOUT(15) => R1IN_1_BCOUT(15),
  BCOUT(16) => R1IN_1_BCOUT(16),
  BCOUT(17) => R1IN_1_BCOUT(17),
  P(0) => PRODUCT(0),
  P(1) => PRODUCT(1),
  P(2) => PRODUCT(2),
  P(3) => PRODUCT(3),
  P(4) => PRODUCT(4),
  P(5) => PRODUCT(5),
  P(6) => PRODUCT(6),
  P(7) => PRODUCT(7),
  P(8) => PRODUCT(8),
  P(9) => PRODUCT(9),
  P(10) => PRODUCT(10),
  P(11) => PRODUCT(11),
  P(12) => PRODUCT(12),
  P(13) => PRODUCT(13),
  P(14) => PRODUCT(14),
  P(15) => PRODUCT(15),
  P(16) => PRODUCT(16),
  P(17) => R1IN_ADD_2,
  P(18) => R1IN_1FF(18),
  P(19) => R1IN_1FF(19),
  P(20) => R1IN_1FF(20),
  P(21) => R1IN_1FF(21),
  P(22) => R1IN_1FF(22),
  P(23) => R1IN_1FF(23),
  P(24) => R1IN_1FF(24),
  P(25) => R1IN_1FF(25),
  P(26) => R1IN_1FF(26),
  P(27) => R1IN_1FF(27),
  P(28) => R1IN_1FF(28),
  P(29) => R1IN_1FF(29),
  P(30) => R1IN_1FF(30),
  P(31) => R1IN_1FF(31),
  P(32) => R1IN_1FF(32),
  P(33) => R1IN_1FF(33),
  P(34) => UC_180,
  P(35) => UC_181,
  P(36) => UC_182,
  P(37) => UC_183,
  P(38) => UC_184,
  P(39) => UC_185,
  P(40) => UC_186,
  P(41) => UC_187,
  P(42) => UC_188,
  P(43) => UC_189,
  P(44) => UC_190,
  P(45) => UC_191,
  P(46) => UC_192,
  P(47) => UC_193,
  PCOUT(0) => R1IN_1_PCOUT(0),
  PCOUT(1) => R1IN_1_PCOUT(1),
  PCOUT(2) => R1IN_1_PCOUT(2),
  PCOUT(3) => R1IN_1_PCOUT(3),
  PCOUT(4) => R1IN_1_PCOUT(4),
  PCOUT(5) => R1IN_1_PCOUT(5),
  PCOUT(6) => R1IN_1_PCOUT(6),
  PCOUT(7) => R1IN_1_PCOUT(7),
  PCOUT(8) => R1IN_1_PCOUT(8),
  PCOUT(9) => R1IN_1_PCOUT(9),
  PCOUT(10) => R1IN_1_PCOUT(10),
  PCOUT(11) => R1IN_1_PCOUT(11),
  PCOUT(12) => R1IN_1_PCOUT(12),
  PCOUT(13) => R1IN_1_PCOUT(13),
  PCOUT(14) => R1IN_1_PCOUT(14),
  PCOUT(15) => R1IN_1_PCOUT(15),
  PCOUT(16) => R1IN_1_PCOUT(16),
  PCOUT(17) => R1IN_1_PCOUT(17),
  PCOUT(18) => R1IN_1_PCOUT(18),
  PCOUT(19) => R1IN_1_PCOUT(19),
  PCOUT(20) => R1IN_1_PCOUT(20),
  PCOUT(21) => R1IN_1_PCOUT(21),
  PCOUT(22) => R1IN_1_PCOUT(22),
  PCOUT(23) => R1IN_1_PCOUT(23),
  PCOUT(24) => R1IN_1_PCOUT(24),
  PCOUT(25) => R1IN_1_PCOUT(25),
  PCOUT(26) => R1IN_1_PCOUT(26),
  PCOUT(27) => R1IN_1_PCOUT(27),
  PCOUT(28) => R1IN_1_PCOUT(28),
  PCOUT(29) => R1IN_1_PCOUT(29),
  PCOUT(30) => R1IN_1_PCOUT(30),
  PCOUT(31) => R1IN_1_PCOUT(31),
  PCOUT(32) => R1IN_1_PCOUT(32),
  PCOUT(33) => R1IN_1_PCOUT(33),
  PCOUT(34) => R1IN_1_PCOUT(34),
  PCOUT(35) => R1IN_1_PCOUT(35),
  PCOUT(36) => R1IN_1_PCOUT(36),
  PCOUT(37) => R1IN_1_PCOUT(37),
  PCOUT(38) => R1IN_1_PCOUT(38),
  PCOUT(39) => R1IN_1_PCOUT(39),
  PCOUT(40) => R1IN_1_PCOUT(40),
  PCOUT(41) => R1IN_1_PCOUT(41),
  PCOUT(42) => R1IN_1_PCOUT(42),
  PCOUT(43) => R1IN_1_PCOUT(43),
  PCOUT(44) => R1IN_1_PCOUT(44),
  PCOUT(45) => R1IN_1_PCOUT(45),
  PCOUT(46) => R1IN_1_PCOUT(46),
  PCOUT(47) => R1IN_1_PCOUT(47));
R1IN_4_3_1q330w: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 0,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => B(34),
  A(1) => B(35),
  A(2) => B(36),
  A(3) => B(37),
  A(4) => B(38),
  A(5) => B(39),
  A(6) => B(40),
  A(7) => B(41),
  A(8) => B(42),
  A(9) => B(43),
  A(10) => B(44),
  A(11) => B(45),
  A(12) => B(46),
  A(13) => B(47),
  A(14) => B(48),
  A(15) => B(49),
  A(16) => B(50),
  A(17) => NN_1,
  B(0) => A(17),
  B(1) => A(18),
  B(2) => A(19),
  B(3) => A(20),
  B(4) => A(21),
  B(5) => A(22),
  B(6) => A(23),
  B(7) => A(24),
  B(8) => A(25),
  B(9) => A(26),
  B(10) => A(27),
  B(11) => A(28),
  B(12) => A(29),
  B(13) => A(30),
  B(14) => A(31),
  B(15) => A(32),
  B(16) => A(33),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => NN_1,
  PCIN(1) => NN_1,
  PCIN(2) => NN_1,
  PCIN(3) => NN_1,
  PCIN(4) => NN_1,
  PCIN(5) => NN_1,
  PCIN(6) => NN_1,
  PCIN(7) => NN_1,
  PCIN(8) => NN_1,
  PCIN(9) => NN_1,
  PCIN(10) => NN_1,
  PCIN(11) => NN_1,
  PCIN(12) => NN_1,
  PCIN(13) => NN_1,
  PCIN(14) => NN_1,
  PCIN(15) => NN_1,
  PCIN(16) => NN_1,
  PCIN(17) => NN_1,
  PCIN(18) => NN_1,
  PCIN(19) => NN_1,
  PCIN(20) => NN_1,
  PCIN(21) => NN_1,
  PCIN(22) => NN_1,
  PCIN(23) => NN_1,
  PCIN(24) => NN_1,
  PCIN(25) => NN_1,
  PCIN(26) => NN_1,
  PCIN(27) => NN_1,
  PCIN(28) => NN_1,
  PCIN(29) => NN_1,
  PCIN(30) => NN_1,
  PCIN(31) => NN_1,
  PCIN(32) => NN_1,
  PCIN(33) => NN_1,
  PCIN(34) => NN_1,
  PCIN(35) => NN_1,
  PCIN(36) => NN_1,
  PCIN(37) => NN_1,
  PCIN(38) => NN_1,
  PCIN(39) => NN_1,
  PCIN(40) => NN_1,
  PCIN(41) => NN_1,
  PCIN(42) => NN_1,
  PCIN(43) => NN_1,
  PCIN(44) => NN_1,
  PCIN(45) => NN_1,
  PCIN(46) => NN_1,
  PCIN(47) => NN_1,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_1,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => NN_1,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => NN_1,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_4_3_1_BCOUT(0),
  BCOUT(1) => R1IN_4_3_1_BCOUT(1),
  BCOUT(2) => R1IN_4_3_1_BCOUT(2),
  BCOUT(3) => R1IN_4_3_1_BCOUT(3),
  BCOUT(4) => R1IN_4_3_1_BCOUT(4),
  BCOUT(5) => R1IN_4_3_1_BCOUT(5),
  BCOUT(6) => R1IN_4_3_1_BCOUT(6),
  BCOUT(7) => R1IN_4_3_1_BCOUT(7),
  BCOUT(8) => R1IN_4_3_1_BCOUT(8),
  BCOUT(9) => R1IN_4_3_1_BCOUT(9),
  BCOUT(10) => R1IN_4_3_1_BCOUT(10),
  BCOUT(11) => R1IN_4_3_1_BCOUT(11),
  BCOUT(12) => R1IN_4_3_1_BCOUT(12),
  BCOUT(13) => R1IN_4_3_1_BCOUT(13),
  BCOUT(14) => R1IN_4_3_1_BCOUT(14),
  BCOUT(15) => R1IN_4_3_1_BCOUT(15),
  BCOUT(16) => R1IN_4_3_1_BCOUT(16),
  BCOUT(17) => R1IN_4_3_1_BCOUT(17),
  P(0) => R1IN_4_3(0),
  P(1) => R1IN_4_3(1),
  P(2) => R1IN_4_3(2),
  P(3) => R1IN_4_3(3),
  P(4) => R1IN_4_3(4),
  P(5) => R1IN_4_3(5),
  P(6) => R1IN_4_3(6),
  P(7) => R1IN_4_3(7),
  P(8) => R1IN_4_3(8),
  P(9) => R1IN_4_3(9),
  P(10) => R1IN_4_3(10),
  P(11) => R1IN_4_3(11),
  P(12) => R1IN_4_3(12),
  P(13) => R1IN_4_3(13),
  P(14) => R1IN_4_3(14),
  P(15) => R1IN_4_3(15),
  P(16) => R1IN_4_3(16),
  P(17) => R1IN_4_3_1(17),
  P(18) => R1IN_4_3_1(18),
  P(19) => R1IN_4_3_1(19),
  P(20) => R1IN_4_3_1(20),
  P(21) => R1IN_4_3_1(21),
  P(22) => R1IN_4_3_1(22),
  P(23) => R1IN_4_3_1(23),
  P(24) => R1IN_4_3_1(24),
  P(25) => R1IN_4_3_1(25),
  P(26) => R1IN_4_3_1(26),
  P(27) => R1IN_4_3_1(27),
  P(28) => R1IN_4_3_1(28),
  P(29) => R1IN_4_3_1(29),
  P(30) => R1IN_4_3_1(30),
  P(31) => R1IN_4_3_1(31),
  P(32) => R1IN_4_3_1(32),
  P(33) => R1IN_4_3_1(33),
  P(34) => UC_166,
  P(35) => UC_167,
  P(36) => UC_168,
  P(37) => UC_169,
  P(38) => UC_170,
  P(39) => UC_171,
  P(40) => UC_172,
  P(41) => UC_173,
  P(42) => UC_174,
  P(43) => UC_175,
  P(44) => UC_176,
  P(45) => UC_177,
  P(46) => UC_178,
  P(47) => UC_179,
  PCOUT(0) => R1IN_4_3_0(0),
  PCOUT(1) => R1IN_4_3_0(1),
  PCOUT(2) => R1IN_4_3_0(2),
  PCOUT(3) => R1IN_4_3_0(3),
  PCOUT(4) => R1IN_4_3_0(4),
  PCOUT(5) => R1IN_4_3_0(5),
  PCOUT(6) => R1IN_4_3_0(6),
  PCOUT(7) => R1IN_4_3_0(7),
  PCOUT(8) => R1IN_4_3_0(8),
  PCOUT(9) => R1IN_4_3_0(9),
  PCOUT(10) => R1IN_4_3_0(10),
  PCOUT(11) => R1IN_4_3_0(11),
  PCOUT(12) => R1IN_4_3_0(12),
  PCOUT(13) => R1IN_4_3_0(13),
  PCOUT(14) => R1IN_4_3_0(14),
  PCOUT(15) => R1IN_4_3_0(15),
  PCOUT(16) => R1IN_4_3_0(16),
  PCOUT(17) => R1IN_4_3_1_0(17),
  PCOUT(18) => R1IN_4_3_1_0(18),
  PCOUT(19) => R1IN_4_3_1_0(19),
  PCOUT(20) => R1IN_4_3_1_0(20),
  PCOUT(21) => R1IN_4_3_1_0(21),
  PCOUT(22) => R1IN_4_3_1_0(22),
  PCOUT(23) => R1IN_4_3_1_0(23),
  PCOUT(24) => R1IN_4_3_1_0(24),
  PCOUT(25) => R1IN_4_3_1_0(25),
  PCOUT(26) => R1IN_4_3_1_0(26),
  PCOUT(27) => R1IN_4_3_1_0(27),
  PCOUT(28) => R1IN_4_3_1_0(28),
  PCOUT(29) => R1IN_4_3_1_0(29),
  PCOUT(30) => R1IN_4_3_1_0(30),
  PCOUT(31) => R1IN_4_3_1_0(31),
  PCOUT(32) => R1IN_4_3_1_0(32),
  PCOUT(33) => R1IN_4_3_1_0(33),
  PCOUT(34) => UC_166_0,
  PCOUT(35) => UC_167_0,
  PCOUT(36) => UC_168_0,
  PCOUT(37) => UC_169_0,
  PCOUT(38) => UC_170_0,
  PCOUT(39) => UC_171_0,
  PCOUT(40) => UC_172_0,
  PCOUT(41) => UC_173_0,
  PCOUT(42) => UC_174_0,
  PCOUT(43) => UC_175_0,
  PCOUT(44) => UC_176_0,
  PCOUT(45) => UC_177_0,
  PCOUT(46) => UC_178_0,
  PCOUT(47) => UC_179_0);
R1IN_4_2_1q330w: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 0,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => A(34),
  A(1) => A(35),
  A(2) => A(36),
  A(3) => A(37),
  A(4) => A(38),
  A(5) => A(39),
  A(6) => A(40),
  A(7) => A(41),
  A(8) => A(42),
  A(9) => A(43),
  A(10) => A(44),
  A(11) => A(45),
  A(12) => A(46),
  A(13) => A(47),
  A(14) => A(48),
  A(15) => A(49),
  A(16) => A(50),
  A(17) => NN_1,
  B(0) => B(17),
  B(1) => B(18),
  B(2) => B(19),
  B(3) => B(20),
  B(4) => B(21),
  B(5) => B(22),
  B(6) => B(23),
  B(7) => B(24),
  B(8) => B(25),
  B(9) => B(26),
  B(10) => B(27),
  B(11) => B(28),
  B(12) => B(29),
  B(13) => B(30),
  B(14) => B(31),
  B(15) => B(32),
  B(16) => B(33),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => NN_1,
  PCIN(1) => NN_1,
  PCIN(2) => NN_1,
  PCIN(3) => NN_1,
  PCIN(4) => NN_1,
  PCIN(5) => NN_1,
  PCIN(6) => NN_1,
  PCIN(7) => NN_1,
  PCIN(8) => NN_1,
  PCIN(9) => NN_1,
  PCIN(10) => NN_1,
  PCIN(11) => NN_1,
  PCIN(12) => NN_1,
  PCIN(13) => NN_1,
  PCIN(14) => NN_1,
  PCIN(15) => NN_1,
  PCIN(16) => NN_1,
  PCIN(17) => NN_1,
  PCIN(18) => NN_1,
  PCIN(19) => NN_1,
  PCIN(20) => NN_1,
  PCIN(21) => NN_1,
  PCIN(22) => NN_1,
  PCIN(23) => NN_1,
  PCIN(24) => NN_1,
  PCIN(25) => NN_1,
  PCIN(26) => NN_1,
  PCIN(27) => NN_1,
  PCIN(28) => NN_1,
  PCIN(29) => NN_1,
  PCIN(30) => NN_1,
  PCIN(31) => NN_1,
  PCIN(32) => NN_1,
  PCIN(33) => NN_1,
  PCIN(34) => NN_1,
  PCIN(35) => NN_1,
  PCIN(36) => NN_1,
  PCIN(37) => NN_1,
  PCIN(38) => NN_1,
  PCIN(39) => NN_1,
  PCIN(40) => NN_1,
  PCIN(41) => NN_1,
  PCIN(42) => NN_1,
  PCIN(43) => NN_1,
  PCIN(44) => NN_1,
  PCIN(45) => NN_1,
  PCIN(46) => NN_1,
  PCIN(47) => NN_1,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_1,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => NN_1,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => NN_1,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_4_2_1_BCOUT(0),
  BCOUT(1) => R1IN_4_2_1_BCOUT(1),
  BCOUT(2) => R1IN_4_2_1_BCOUT(2),
  BCOUT(3) => R1IN_4_2_1_BCOUT(3),
  BCOUT(4) => R1IN_4_2_1_BCOUT(4),
  BCOUT(5) => R1IN_4_2_1_BCOUT(5),
  BCOUT(6) => R1IN_4_2_1_BCOUT(6),
  BCOUT(7) => R1IN_4_2_1_BCOUT(7),
  BCOUT(8) => R1IN_4_2_1_BCOUT(8),
  BCOUT(9) => R1IN_4_2_1_BCOUT(9),
  BCOUT(10) => R1IN_4_2_1_BCOUT(10),
  BCOUT(11) => R1IN_4_2_1_BCOUT(11),
  BCOUT(12) => R1IN_4_2_1_BCOUT(12),
  BCOUT(13) => R1IN_4_2_1_BCOUT(13),
  BCOUT(14) => R1IN_4_2_1_BCOUT(14),
  BCOUT(15) => R1IN_4_2_1_BCOUT(15),
  BCOUT(16) => R1IN_4_2_1_BCOUT(16),
  BCOUT(17) => R1IN_4_2_1_BCOUT(17),
  P(0) => R1IN_4_2(0),
  P(1) => R1IN_4_2(1),
  P(2) => R1IN_4_2(2),
  P(3) => R1IN_4_2(3),
  P(4) => R1IN_4_2(4),
  P(5) => R1IN_4_2(5),
  P(6) => R1IN_4_2(6),
  P(7) => R1IN_4_2(7),
  P(8) => R1IN_4_2(8),
  P(9) => R1IN_4_2(9),
  P(10) => R1IN_4_2(10),
  P(11) => R1IN_4_2(11),
  P(12) => R1IN_4_2(12),
  P(13) => R1IN_4_2(13),
  P(14) => R1IN_4_2(14),
  P(15) => R1IN_4_2(15),
  P(16) => R1IN_4_2(16),
  P(17) => R1IN_4_2_1(17),
  P(18) => R1IN_4_2_1(18),
  P(19) => R1IN_4_2_1(19),
  P(20) => R1IN_4_2_1(20),
  P(21) => R1IN_4_2_1(21),
  P(22) => R1IN_4_2_1(22),
  P(23) => R1IN_4_2_1(23),
  P(24) => R1IN_4_2_1(24),
  P(25) => R1IN_4_2_1(25),
  P(26) => R1IN_4_2_1(26),
  P(27) => R1IN_4_2_1(27),
  P(28) => R1IN_4_2_1(28),
  P(29) => R1IN_4_2_1(29),
  P(30) => R1IN_4_2_1(30),
  P(31) => R1IN_4_2_1(31),
  P(32) => R1IN_4_2_1(32),
  P(33) => R1IN_4_2_1(33),
  P(34) => UC_152,
  P(35) => UC_153,
  P(36) => UC_154,
  P(37) => UC_155,
  P(38) => UC_156,
  P(39) => UC_157,
  P(40) => UC_158,
  P(41) => UC_159,
  P(42) => UC_160,
  P(43) => UC_161,
  P(44) => UC_162,
  P(45) => UC_163,
  P(46) => UC_164,
  P(47) => UC_165,
  PCOUT(0) => R1IN_4_2_0(0),
  PCOUT(1) => R1IN_4_2_0(1),
  PCOUT(2) => R1IN_4_2_0(2),
  PCOUT(3) => R1IN_4_2_0(3),
  PCOUT(4) => R1IN_4_2_0(4),
  PCOUT(5) => R1IN_4_2_0(5),
  PCOUT(6) => R1IN_4_2_0(6),
  PCOUT(7) => R1IN_4_2_0(7),
  PCOUT(8) => R1IN_4_2_0(8),
  PCOUT(9) => R1IN_4_2_0(9),
  PCOUT(10) => R1IN_4_2_0(10),
  PCOUT(11) => R1IN_4_2_0(11),
  PCOUT(12) => R1IN_4_2_0(12),
  PCOUT(13) => R1IN_4_2_0(13),
  PCOUT(14) => R1IN_4_2_0(14),
  PCOUT(15) => R1IN_4_2_0(15),
  PCOUT(16) => R1IN_4_2_0(16),
  PCOUT(17) => R1IN_4_2_1_0(17),
  PCOUT(18) => R1IN_4_2_1_0(18),
  PCOUT(19) => R1IN_4_2_1_0(19),
  PCOUT(20) => R1IN_4_2_1_0(20),
  PCOUT(21) => R1IN_4_2_1_0(21),
  PCOUT(22) => R1IN_4_2_1_0(22),
  PCOUT(23) => R1IN_4_2_1_0(23),
  PCOUT(24) => R1IN_4_2_1_0(24),
  PCOUT(25) => R1IN_4_2_1_0(25),
  PCOUT(26) => R1IN_4_2_1_0(26),
  PCOUT(27) => R1IN_4_2_1_0(27),
  PCOUT(28) => R1IN_4_2_1_0(28),
  PCOUT(29) => R1IN_4_2_1_0(29),
  PCOUT(30) => R1IN_4_2_1_0(30),
  PCOUT(31) => R1IN_4_2_1_0(31),
  PCOUT(32) => R1IN_4_2_1_0(32),
  PCOUT(33) => R1IN_4_2_1_0(33),
  PCOUT(34) => UC_152_0,
  PCOUT(35) => UC_153_0,
  PCOUT(36) => UC_154_0,
  PCOUT(37) => UC_155_0,
  PCOUT(38) => UC_156_0,
  PCOUT(39) => UC_157_0,
  PCOUT(40) => UC_158_0,
  PCOUT(41) => UC_159_0,
  PCOUT(42) => UC_160_0,
  PCOUT(43) => UC_161_0,
  PCOUT(44) => UC_162_0,
  PCOUT(45) => UC_163_0,
  PCOUT(46) => UC_164_0,
  PCOUT(47) => UC_165_0);
R1IN_3_2_1q330w: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 0,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => B(34),
  A(1) => B(35),
  A(2) => B(36),
  A(3) => B(37),
  A(4) => B(38),
  A(5) => B(39),
  A(6) => B(40),
  A(7) => B(41),
  A(8) => B(42),
  A(9) => B(43),
  A(10) => B(44),
  A(11) => B(45),
  A(12) => B(46),
  A(13) => B(47),
  A(14) => B(48),
  A(15) => B(49),
  A(16) => B(50),
  A(17) => NN_1,
  B(0) => A(0),
  B(1) => A(1),
  B(2) => A(2),
  B(3) => A(3),
  B(4) => A(4),
  B(5) => A(5),
  B(6) => A(6),
  B(7) => A(7),
  B(8) => A(8),
  B(9) => A(9),
  B(10) => A(10),
  B(11) => A(11),
  B(12) => A(12),
  B(13) => A(13),
  B(14) => A(14),
  B(15) => A(15),
  B(16) => A(16),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => NN_1,
  PCIN(1) => NN_1,
  PCIN(2) => NN_1,
  PCIN(3) => NN_1,
  PCIN(4) => NN_1,
  PCIN(5) => NN_1,
  PCIN(6) => NN_1,
  PCIN(7) => NN_1,
  PCIN(8) => NN_1,
  PCIN(9) => NN_1,
  PCIN(10) => NN_1,
  PCIN(11) => NN_1,
  PCIN(12) => NN_1,
  PCIN(13) => NN_1,
  PCIN(14) => NN_1,
  PCIN(15) => NN_1,
  PCIN(16) => NN_1,
  PCIN(17) => NN_1,
  PCIN(18) => NN_1,
  PCIN(19) => NN_1,
  PCIN(20) => NN_1,
  PCIN(21) => NN_1,
  PCIN(22) => NN_1,
  PCIN(23) => NN_1,
  PCIN(24) => NN_1,
  PCIN(25) => NN_1,
  PCIN(26) => NN_1,
  PCIN(27) => NN_1,
  PCIN(28) => NN_1,
  PCIN(29) => NN_1,
  PCIN(30) => NN_1,
  PCIN(31) => NN_1,
  PCIN(32) => NN_1,
  PCIN(33) => NN_1,
  PCIN(34) => NN_1,
  PCIN(35) => NN_1,
  PCIN(36) => NN_1,
  PCIN(37) => NN_1,
  PCIN(38) => NN_1,
  PCIN(39) => NN_1,
  PCIN(40) => NN_1,
  PCIN(41) => NN_1,
  PCIN(42) => NN_1,
  PCIN(43) => NN_1,
  PCIN(44) => NN_1,
  PCIN(45) => NN_1,
  PCIN(46) => NN_1,
  PCIN(47) => NN_1,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_1,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => NN_1,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => NN_1,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_3_2_1_BCOUT(0),
  BCOUT(1) => R1IN_3_2_1_BCOUT(1),
  BCOUT(2) => R1IN_3_2_1_BCOUT(2),
  BCOUT(3) => R1IN_3_2_1_BCOUT(3),
  BCOUT(4) => R1IN_3_2_1_BCOUT(4),
  BCOUT(5) => R1IN_3_2_1_BCOUT(5),
  BCOUT(6) => R1IN_3_2_1_BCOUT(6),
  BCOUT(7) => R1IN_3_2_1_BCOUT(7),
  BCOUT(8) => R1IN_3_2_1_BCOUT(8),
  BCOUT(9) => R1IN_3_2_1_BCOUT(9),
  BCOUT(10) => R1IN_3_2_1_BCOUT(10),
  BCOUT(11) => R1IN_3_2_1_BCOUT(11),
  BCOUT(12) => R1IN_3_2_1_BCOUT(12),
  BCOUT(13) => R1IN_3_2_1_BCOUT(13),
  BCOUT(14) => R1IN_3_2_1_BCOUT(14),
  BCOUT(15) => R1IN_3_2_1_BCOUT(15),
  BCOUT(16) => R1IN_3_2_1_BCOUT(16),
  BCOUT(17) => R1IN_3_2_1_BCOUT(17),
  P(0) => R1IN_3_2(0),
  P(1) => R1IN_3_2(1),
  P(2) => R1IN_3_2(2),
  P(3) => R1IN_3_2(3),
  P(4) => R1IN_3_2(4),
  P(5) => R1IN_3_2(5),
  P(6) => R1IN_3_2(6),
  P(7) => R1IN_3_2(7),
  P(8) => R1IN_3_2(8),
  P(9) => R1IN_3_2(9),
  P(10) => R1IN_3_2(10),
  P(11) => R1IN_3_2(11),
  P(12) => R1IN_3_2(12),
  P(13) => R1IN_3_2(13),
  P(14) => R1IN_3_2(14),
  P(15) => R1IN_3_2(15),
  P(16) => R1IN_3_2(16),
  P(17) => R1IN_3_2_1(17),
  P(18) => R1IN_3_2_1(18),
  P(19) => R1IN_3_2_1(19),
  P(20) => R1IN_3_2_1(20),
  P(21) => R1IN_3_2_1(21),
  P(22) => R1IN_3_2_1(22),
  P(23) => R1IN_3_2_1(23),
  P(24) => R1IN_3_2_1(24),
  P(25) => R1IN_3_2_1(25),
  P(26) => R1IN_3_2_1(26),
  P(27) => R1IN_3_2_1(27),
  P(28) => R1IN_3_2_1(28),
  P(29) => R1IN_3_2_1(29),
  P(30) => R1IN_3_2_1(30),
  P(31) => R1IN_3_2_1(31),
  P(32) => R1IN_3_2_1(32),
  P(33) => R1IN_3_2_1(33),
  P(34) => UC_138,
  P(35) => UC_139,
  P(36) => UC_140,
  P(37) => UC_141,
  P(38) => UC_142,
  P(39) => UC_143,
  P(40) => UC_144,
  P(41) => UC_145,
  P(42) => UC_146,
  P(43) => UC_147,
  P(44) => UC_148,
  P(45) => UC_149,
  P(46) => UC_150,
  P(47) => UC_151,
  PCOUT(0) => R1IN_3_2_0(0),
  PCOUT(1) => R1IN_3_2_0(1),
  PCOUT(2) => R1IN_3_2_0(2),
  PCOUT(3) => R1IN_3_2_0(3),
  PCOUT(4) => R1IN_3_2_0(4),
  PCOUT(5) => R1IN_3_2_0(5),
  PCOUT(6) => R1IN_3_2_0(6),
  PCOUT(7) => R1IN_3_2_0(7),
  PCOUT(8) => R1IN_3_2_0(8),
  PCOUT(9) => R1IN_3_2_0(9),
  PCOUT(10) => R1IN_3_2_0(10),
  PCOUT(11) => R1IN_3_2_0(11),
  PCOUT(12) => R1IN_3_2_0(12),
  PCOUT(13) => R1IN_3_2_0(13),
  PCOUT(14) => R1IN_3_2_0(14),
  PCOUT(15) => R1IN_3_2_0(15),
  PCOUT(16) => R1IN_3_2_0(16),
  PCOUT(17) => R1IN_3_2_1_0(17),
  PCOUT(18) => R1IN_3_2_1_0(18),
  PCOUT(19) => R1IN_3_2_1_0(19),
  PCOUT(20) => R1IN_3_2_1_0(20),
  PCOUT(21) => R1IN_3_2_1_0(21),
  PCOUT(22) => R1IN_3_2_1_0(22),
  PCOUT(23) => R1IN_3_2_1_0(23),
  PCOUT(24) => R1IN_3_2_1_0(24),
  PCOUT(25) => R1IN_3_2_1_0(25),
  PCOUT(26) => R1IN_3_2_1_0(26),
  PCOUT(27) => R1IN_3_2_1_0(27),
  PCOUT(28) => R1IN_3_2_1_0(28),
  PCOUT(29) => R1IN_3_2_1_0(29),
  PCOUT(30) => R1IN_3_2_1_0(30),
  PCOUT(31) => R1IN_3_2_1_0(31),
  PCOUT(32) => R1IN_3_2_1_0(32),
  PCOUT(33) => R1IN_3_2_1_0(33),
  PCOUT(34) => UC_138_0,
  PCOUT(35) => UC_139_0,
  PCOUT(36) => UC_140_0,
  PCOUT(37) => UC_141_0,
  PCOUT(38) => UC_142_0,
  PCOUT(39) => UC_143_0,
  PCOUT(40) => UC_144_0,
  PCOUT(41) => UC_145_0,
  PCOUT(42) => UC_146_0,
  PCOUT(43) => UC_147_0,
  PCOUT(44) => UC_148_0,
  PCOUT(45) => UC_149_0,
  PCOUT(46) => UC_150_0,
  PCOUT(47) => UC_151_0);
R1IN_2_2_1q330w: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 0,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => A(34),
  A(1) => A(35),
  A(2) => A(36),
  A(3) => A(37),
  A(4) => A(38),
  A(5) => A(39),
  A(6) => A(40),
  A(7) => A(41),
  A(8) => A(42),
  A(9) => A(43),
  A(10) => A(44),
  A(11) => A(45),
  A(12) => A(46),
  A(13) => A(47),
  A(14) => A(48),
  A(15) => A(49),
  A(16) => A(50),
  A(17) => NN_1,
  B(0) => B(0),
  B(1) => B(1),
  B(2) => B(2),
  B(3) => B(3),
  B(4) => B(4),
  B(5) => B(5),
  B(6) => B(6),
  B(7) => B(7),
  B(8) => B(8),
  B(9) => B(9),
  B(10) => B(10),
  B(11) => B(11),
  B(12) => B(12),
  B(13) => B(13),
  B(14) => B(14),
  B(15) => B(15),
  B(16) => B(16),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => NN_1,
  PCIN(1) => NN_1,
  PCIN(2) => NN_1,
  PCIN(3) => NN_1,
  PCIN(4) => NN_1,
  PCIN(5) => NN_1,
  PCIN(6) => NN_1,
  PCIN(7) => NN_1,
  PCIN(8) => NN_1,
  PCIN(9) => NN_1,
  PCIN(10) => NN_1,
  PCIN(11) => NN_1,
  PCIN(12) => NN_1,
  PCIN(13) => NN_1,
  PCIN(14) => NN_1,
  PCIN(15) => NN_1,
  PCIN(16) => NN_1,
  PCIN(17) => NN_1,
  PCIN(18) => NN_1,
  PCIN(19) => NN_1,
  PCIN(20) => NN_1,
  PCIN(21) => NN_1,
  PCIN(22) => NN_1,
  PCIN(23) => NN_1,
  PCIN(24) => NN_1,
  PCIN(25) => NN_1,
  PCIN(26) => NN_1,
  PCIN(27) => NN_1,
  PCIN(28) => NN_1,
  PCIN(29) => NN_1,
  PCIN(30) => NN_1,
  PCIN(31) => NN_1,
  PCIN(32) => NN_1,
  PCIN(33) => NN_1,
  PCIN(34) => NN_1,
  PCIN(35) => NN_1,
  PCIN(36) => NN_1,
  PCIN(37) => NN_1,
  PCIN(38) => NN_1,
  PCIN(39) => NN_1,
  PCIN(40) => NN_1,
  PCIN(41) => NN_1,
  PCIN(42) => NN_1,
  PCIN(43) => NN_1,
  PCIN(44) => NN_1,
  PCIN(45) => NN_1,
  PCIN(46) => NN_1,
  PCIN(47) => NN_1,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_1,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => NN_1,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => NN_1,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_2_2_1_BCOUT(0),
  BCOUT(1) => R1IN_2_2_1_BCOUT(1),
  BCOUT(2) => R1IN_2_2_1_BCOUT(2),
  BCOUT(3) => R1IN_2_2_1_BCOUT(3),
  BCOUT(4) => R1IN_2_2_1_BCOUT(4),
  BCOUT(5) => R1IN_2_2_1_BCOUT(5),
  BCOUT(6) => R1IN_2_2_1_BCOUT(6),
  BCOUT(7) => R1IN_2_2_1_BCOUT(7),
  BCOUT(8) => R1IN_2_2_1_BCOUT(8),
  BCOUT(9) => R1IN_2_2_1_BCOUT(9),
  BCOUT(10) => R1IN_2_2_1_BCOUT(10),
  BCOUT(11) => R1IN_2_2_1_BCOUT(11),
  BCOUT(12) => R1IN_2_2_1_BCOUT(12),
  BCOUT(13) => R1IN_2_2_1_BCOUT(13),
  BCOUT(14) => R1IN_2_2_1_BCOUT(14),
  BCOUT(15) => R1IN_2_2_1_BCOUT(15),
  BCOUT(16) => R1IN_2_2_1_BCOUT(16),
  BCOUT(17) => R1IN_2_2_1_BCOUT(17),
  P(0) => R1IN_2_2(0),
  P(1) => R1IN_2_2(1),
  P(2) => R1IN_2_2(2),
  P(3) => R1IN_2_2(3),
  P(4) => R1IN_2_2(4),
  P(5) => R1IN_2_2(5),
  P(6) => R1IN_2_2(6),
  P(7) => R1IN_2_2(7),
  P(8) => R1IN_2_2(8),
  P(9) => R1IN_2_2(9),
  P(10) => R1IN_2_2(10),
  P(11) => R1IN_2_2(11),
  P(12) => R1IN_2_2(12),
  P(13) => R1IN_2_2(13),
  P(14) => R1IN_2_2(14),
  P(15) => R1IN_2_2(15),
  P(16) => R1IN_2_2(16),
  P(17) => R1IN_2_2_1(17),
  P(18) => R1IN_2_2_1(18),
  P(19) => R1IN_2_2_1(19),
  P(20) => R1IN_2_2_1(20),
  P(21) => R1IN_2_2_1(21),
  P(22) => R1IN_2_2_1(22),
  P(23) => R1IN_2_2_1(23),
  P(24) => R1IN_2_2_1(24),
  P(25) => R1IN_2_2_1(25),
  P(26) => R1IN_2_2_1(26),
  P(27) => R1IN_2_2_1(27),
  P(28) => R1IN_2_2_1(28),
  P(29) => R1IN_2_2_1(29),
  P(30) => R1IN_2_2_1(30),
  P(31) => R1IN_2_2_1(31),
  P(32) => R1IN_2_2_1(32),
  P(33) => R1IN_2_2_1(33),
  P(34) => UC_124,
  P(35) => UC_125,
  P(36) => UC_126,
  P(37) => UC_127,
  P(38) => UC_128,
  P(39) => UC_129,
  P(40) => UC_130,
  P(41) => UC_131,
  P(42) => UC_132,
  P(43) => UC_133,
  P(44) => UC_134,
  P(45) => UC_135,
  P(46) => UC_136,
  P(47) => UC_137,
  PCOUT(0) => R1IN_2_2_0(0),
  PCOUT(1) => R1IN_2_2_0(1),
  PCOUT(2) => R1IN_2_2_0(2),
  PCOUT(3) => R1IN_2_2_0(3),
  PCOUT(4) => R1IN_2_2_0(4),
  PCOUT(5) => R1IN_2_2_0(5),
  PCOUT(6) => R1IN_2_2_0(6),
  PCOUT(7) => R1IN_2_2_0(7),
  PCOUT(8) => R1IN_2_2_0(8),
  PCOUT(9) => R1IN_2_2_0(9),
  PCOUT(10) => R1IN_2_2_0(10),
  PCOUT(11) => R1IN_2_2_0(11),
  PCOUT(12) => R1IN_2_2_0(12),
  PCOUT(13) => R1IN_2_2_0(13),
  PCOUT(14) => R1IN_2_2_0(14),
  PCOUT(15) => R1IN_2_2_0(15),
  PCOUT(16) => R1IN_2_2_0(16),
  PCOUT(17) => R1IN_2_2_1_0(17),
  PCOUT(18) => R1IN_2_2_1_0(18),
  PCOUT(19) => R1IN_2_2_1_0(19),
  PCOUT(20) => R1IN_2_2_1_0(20),
  PCOUT(21) => R1IN_2_2_1_0(21),
  PCOUT(22) => R1IN_2_2_1_0(22),
  PCOUT(23) => R1IN_2_2_1_0(23),
  PCOUT(24) => R1IN_2_2_1_0(24),
  PCOUT(25) => R1IN_2_2_1_0(25),
  PCOUT(26) => R1IN_2_2_1_0(26),
  PCOUT(27) => R1IN_2_2_1_0(27),
  PCOUT(28) => R1IN_2_2_1_0(28),
  PCOUT(29) => R1IN_2_2_1_0(29),
  PCOUT(30) => R1IN_2_2_1_0(30),
  PCOUT(31) => R1IN_2_2_1_0(31),
  PCOUT(32) => R1IN_2_2_1_0(32),
  PCOUT(33) => R1IN_2_2_1_0(33),
  PCOUT(34) => UC_124_0,
  PCOUT(35) => UC_125_0,
  PCOUT(36) => UC_126_0,
  PCOUT(37) => UC_127_0,
  PCOUT(38) => UC_128_0,
  PCOUT(39) => UC_129_0,
  PCOUT(40) => UC_130_0,
  PCOUT(41) => UC_131_0,
  PCOUT(42) => UC_132_0,
  PCOUT(43) => UC_133_0,
  PCOUT(44) => UC_134_0,
  PCOUT(45) => UC_135_0,
  PCOUT(46) => UC_136_0,
  PCOUT(47) => UC_137_0);
R1IN_4_4_2q260w: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 0,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => A(51),
  A(1) => A(52),
  A(2) => A(53),
  A(3) => A(54),
  A(4) => A(55),
  A(5) => A(56),
  A(6) => A(57),
  A(7) => A(58),
  A(8) => A(59),
  A(9) => A(60),
  A(10) => NN_1,
  A(11) => NN_1,
  A(12) => NN_1,
  A(13) => NN_1,
  A(14) => NN_1,
  A(15) => NN_1,
  A(16) => NN_1,
  A(17) => NN_1,
  B(0) => B(34),
  B(1) => B(35),
  B(2) => B(36),
  B(3) => B(37),
  B(4) => B(38),
  B(5) => B(39),
  B(6) => B(40),
  B(7) => B(41),
  B(8) => B(42),
  B(9) => B(43),
  B(10) => B(44),
  B(11) => B(45),
  B(12) => B(46),
  B(13) => B(47),
  B(14) => B(48),
  B(15) => B(49),
  B(16) => B(50),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => NN_1,
  PCIN(1) => NN_1,
  PCIN(2) => NN_1,
  PCIN(3) => NN_1,
  PCIN(4) => NN_1,
  PCIN(5) => NN_1,
  PCIN(6) => NN_1,
  PCIN(7) => NN_1,
  PCIN(8) => NN_1,
  PCIN(9) => NN_1,
  PCIN(10) => NN_1,
  PCIN(11) => NN_1,
  PCIN(12) => NN_1,
  PCIN(13) => NN_1,
  PCIN(14) => NN_1,
  PCIN(15) => NN_1,
  PCIN(16) => NN_1,
  PCIN(17) => NN_1,
  PCIN(18) => NN_1,
  PCIN(19) => NN_1,
  PCIN(20) => NN_1,
  PCIN(21) => NN_1,
  PCIN(22) => NN_1,
  PCIN(23) => NN_1,
  PCIN(24) => NN_1,
  PCIN(25) => NN_1,
  PCIN(26) => NN_1,
  PCIN(27) => NN_1,
  PCIN(28) => NN_1,
  PCIN(29) => NN_1,
  PCIN(30) => NN_1,
  PCIN(31) => NN_1,
  PCIN(32) => NN_1,
  PCIN(33) => NN_1,
  PCIN(34) => NN_1,
  PCIN(35) => NN_1,
  PCIN(36) => NN_1,
  PCIN(37) => NN_1,
  PCIN(38) => NN_1,
  PCIN(39) => NN_1,
  PCIN(40) => NN_1,
  PCIN(41) => NN_1,
  PCIN(42) => NN_1,
  PCIN(43) => NN_1,
  PCIN(44) => NN_1,
  PCIN(45) => NN_1,
  PCIN(46) => NN_1,
  PCIN(47) => NN_1,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_1,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => NN_1,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => NN_1,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_4_4_2_BCOUT(0),
  BCOUT(1) => R1IN_4_4_2_BCOUT(1),
  BCOUT(2) => R1IN_4_4_2_BCOUT(2),
  BCOUT(3) => R1IN_4_4_2_BCOUT(3),
  BCOUT(4) => R1IN_4_4_2_BCOUT(4),
  BCOUT(5) => R1IN_4_4_2_BCOUT(5),
  BCOUT(6) => R1IN_4_4_2_BCOUT(6),
  BCOUT(7) => R1IN_4_4_2_BCOUT(7),
  BCOUT(8) => R1IN_4_4_2_BCOUT(8),
  BCOUT(9) => R1IN_4_4_2_BCOUT(9),
  BCOUT(10) => R1IN_4_4_2_BCOUT(10),
  BCOUT(11) => R1IN_4_4_2_BCOUT(11),
  BCOUT(12) => R1IN_4_4_2_BCOUT(12),
  BCOUT(13) => R1IN_4_4_2_BCOUT(13),
  BCOUT(14) => R1IN_4_4_2_BCOUT(14),
  BCOUT(15) => R1IN_4_4_2_BCOUT(15),
  BCOUT(16) => R1IN_4_4_2_BCOUT(16),
  BCOUT(17) => R1IN_4_4_2_BCOUT(17),
  P(0) => R1IN_4_4_2(0),
  P(1) => R1IN_4_4_2(1),
  P(2) => R1IN_4_4_2(2),
  P(3) => R1IN_4_4_2(3),
  P(4) => R1IN_4_4_2(4),
  P(5) => R1IN_4_4_2(5),
  P(6) => R1IN_4_4_2(6),
  P(7) => R1IN_4_4_2(7),
  P(8) => R1IN_4_4_2(8),
  P(9) => R1IN_4_4_2(9),
  P(10) => R1IN_4_4_2(10),
  P(11) => R1IN_4_4_2(11),
  P(12) => R1IN_4_4_2(12),
  P(13) => R1IN_4_4_2(13),
  P(14) => R1IN_4_4_2(14),
  P(15) => R1IN_4_4_2(15),
  P(16) => R1IN_4_4_2(16),
  P(17) => R1IN_4_4_2(17),
  P(18) => R1IN_4_4_2(18),
  P(19) => R1IN_4_4_2(19),
  P(20) => R1IN_4_4_2(20),
  P(21) => R1IN_4_4_2(21),
  P(22) => R1IN_4_4_2(22),
  P(23) => R1IN_4_4_2(23),
  P(24) => R1IN_4_4_2(24),
  P(25) => R1IN_4_4_2(25),
  P(26) => R1IN_4_4_2(26),
  P(27) => UC_103,
  P(28) => UC_104,
  P(29) => UC_105,
  P(30) => UC_106,
  P(31) => UC_107,
  P(32) => UC_108,
  P(33) => UC_109,
  P(34) => UC_110,
  P(35) => UC_111,
  P(36) => UC_112,
  P(37) => UC_113,
  P(38) => UC_114,
  P(39) => UC_115,
  P(40) => UC_116,
  P(41) => UC_117,
  P(42) => UC_118,
  P(43) => UC_119,
  P(44) => UC_120,
  P(45) => UC_121,
  P(46) => UC_122,
  P(47) => UC_123,
  PCOUT(0) => R1IN_4_4_2_0(0),
  PCOUT(1) => R1IN_4_4_2_0(1),
  PCOUT(2) => R1IN_4_4_2_0(2),
  PCOUT(3) => R1IN_4_4_2_0(3),
  PCOUT(4) => R1IN_4_4_2_0(4),
  PCOUT(5) => R1IN_4_4_2_0(5),
  PCOUT(6) => R1IN_4_4_2_0(6),
  PCOUT(7) => R1IN_4_4_2_0(7),
  PCOUT(8) => R1IN_4_4_2_0(8),
  PCOUT(9) => R1IN_4_4_2_0(9),
  PCOUT(10) => R1IN_4_4_2_0(10),
  PCOUT(11) => R1IN_4_4_2_0(11),
  PCOUT(12) => R1IN_4_4_2_0(12),
  PCOUT(13) => R1IN_4_4_2_0(13),
  PCOUT(14) => R1IN_4_4_2_0(14),
  PCOUT(15) => R1IN_4_4_2_0(15),
  PCOUT(16) => R1IN_4_4_2_0(16),
  PCOUT(17) => R1IN_4_4_2_0(17),
  PCOUT(18) => R1IN_4_4_2_0(18),
  PCOUT(19) => R1IN_4_4_2_0(19),
  PCOUT(20) => R1IN_4_4_2_0(20),
  PCOUT(21) => R1IN_4_4_2_0(21),
  PCOUT(22) => R1IN_4_4_2_0(22),
  PCOUT(23) => R1IN_4_4_2_0(23),
  PCOUT(24) => R1IN_4_4_2_0(24),
  PCOUT(25) => R1IN_4_4_2_0(25),
  PCOUT(26) => R1IN_4_4_2_0(26),
  PCOUT(27) => UC_103_0,
  PCOUT(28) => UC_104_0,
  PCOUT(29) => UC_105_0,
  PCOUT(30) => UC_106_0,
  PCOUT(31) => UC_107_0,
  PCOUT(32) => UC_108_0,
  PCOUT(33) => UC_109_0,
  PCOUT(34) => UC_110_0,
  PCOUT(35) => UC_111_0,
  PCOUT(36) => UC_112_0,
  PCOUT(37) => UC_113_0,
  PCOUT(38) => UC_114_0,
  PCOUT(39) => UC_115_0,
  PCOUT(40) => UC_116_0,
  PCOUT(41) => UC_117_0,
  PCOUT(42) => UC_118_0,
  PCOUT(43) => UC_119_0,
  PCOUT(44) => UC_120_0,
  PCOUT(45) => UC_121_0,
  PCOUT(46) => UC_122_0,
  PCOUT(47) => UC_123_0);
R1IN_4_3_ADD_1q260w: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 1,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => B(51),
  A(1) => B(52),
  A(2) => B(53),
  A(3) => B(54),
  A(4) => B(55),
  A(5) => B(56),
  A(6) => B(57),
  A(7) => B(58),
  A(8) => B(59),
  A(9) => B(60),
  A(10) => NN_1,
  A(11) => NN_1,
  A(12) => NN_1,
  A(13) => NN_1,
  A(14) => NN_1,
  A(15) => NN_1,
  A(16) => NN_1,
  A(17) => NN_1,
  B(0) => A(17),
  B(1) => A(18),
  B(2) => A(19),
  B(3) => A(20),
  B(4) => A(21),
  B(5) => A(22),
  B(6) => A(23),
  B(7) => A(24),
  B(8) => A(25),
  B(9) => A(26),
  B(10) => A(27),
  B(11) => A(28),
  B(12) => A(29),
  B(13) => A(30),
  B(14) => A(31),
  B(15) => A(32),
  B(16) => A(33),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => R1IN_4_3_0(0),
  PCIN(1) => R1IN_4_3_0(1),
  PCIN(2) => R1IN_4_3_0(2),
  PCIN(3) => R1IN_4_3_0(3),
  PCIN(4) => R1IN_4_3_0(4),
  PCIN(5) => R1IN_4_3_0(5),
  PCIN(6) => R1IN_4_3_0(6),
  PCIN(7) => R1IN_4_3_0(7),
  PCIN(8) => R1IN_4_3_0(8),
  PCIN(9) => R1IN_4_3_0(9),
  PCIN(10) => R1IN_4_3_0(10),
  PCIN(11) => R1IN_4_3_0(11),
  PCIN(12) => R1IN_4_3_0(12),
  PCIN(13) => R1IN_4_3_0(13),
  PCIN(14) => R1IN_4_3_0(14),
  PCIN(15) => R1IN_4_3_0(15),
  PCIN(16) => R1IN_4_3_0(16),
  PCIN(17) => R1IN_4_3_1_0(17),
  PCIN(18) => R1IN_4_3_1_0(18),
  PCIN(19) => R1IN_4_3_1_0(19),
  PCIN(20) => R1IN_4_3_1_0(20),
  PCIN(21) => R1IN_4_3_1_0(21),
  PCIN(22) => R1IN_4_3_1_0(22),
  PCIN(23) => R1IN_4_3_1_0(23),
  PCIN(24) => R1IN_4_3_1_0(24),
  PCIN(25) => R1IN_4_3_1_0(25),
  PCIN(26) => R1IN_4_3_1_0(26),
  PCIN(27) => R1IN_4_3_1_0(27),
  PCIN(28) => R1IN_4_3_1_0(28),
  PCIN(29) => R1IN_4_3_1_0(29),
  PCIN(30) => R1IN_4_3_1_0(30),
  PCIN(31) => R1IN_4_3_1_0(31),
  PCIN(32) => R1IN_4_3_1_0(32),
  PCIN(33) => R1IN_4_3_1_0(33),
  PCIN(34) => UC_166_0,
  PCIN(35) => UC_167_0,
  PCIN(36) => UC_168_0,
  PCIN(37) => UC_169_0,
  PCIN(38) => UC_170_0,
  PCIN(39) => UC_171_0,
  PCIN(40) => UC_172_0,
  PCIN(41) => UC_173_0,
  PCIN(42) => UC_174_0,
  PCIN(43) => UC_175_0,
  PCIN(44) => UC_176_0,
  PCIN(45) => UC_177_0,
  PCIN(46) => UC_178_0,
  PCIN(47) => UC_179_0,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_2,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_2,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => CLK,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => EN,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_4_3_ADD_1_BCOUT(0),
  BCOUT(1) => R1IN_4_3_ADD_1_BCOUT(1),
  BCOUT(2) => R1IN_4_3_ADD_1_BCOUT(2),
  BCOUT(3) => R1IN_4_3_ADD_1_BCOUT(3),
  BCOUT(4) => R1IN_4_3_ADD_1_BCOUT(4),
  BCOUT(5) => R1IN_4_3_ADD_1_BCOUT(5),
  BCOUT(6) => R1IN_4_3_ADD_1_BCOUT(6),
  BCOUT(7) => R1IN_4_3_ADD_1_BCOUT(7),
  BCOUT(8) => R1IN_4_3_ADD_1_BCOUT(8),
  BCOUT(9) => R1IN_4_3_ADD_1_BCOUT(9),
  BCOUT(10) => R1IN_4_3_ADD_1_BCOUT(10),
  BCOUT(11) => R1IN_4_3_ADD_1_BCOUT(11),
  BCOUT(12) => R1IN_4_3_ADD_1_BCOUT(12),
  BCOUT(13) => R1IN_4_3_ADD_1_BCOUT(13),
  BCOUT(14) => R1IN_4_3_ADD_1_BCOUT(14),
  BCOUT(15) => R1IN_4_3_ADD_1_BCOUT(15),
  BCOUT(16) => R1IN_4_3_ADD_1_BCOUT(16),
  BCOUT(17) => R1IN_4_3_ADD_1_BCOUT(17),
  P(0) => R1IN_4_3F(17),
  P(1) => R1IN_4_3F(18),
  P(2) => R1IN_4_3F(19),
  P(3) => R1IN_4_3F(20),
  P(4) => R1IN_4_3F(21),
  P(5) => R1IN_4_3F(22),
  P(6) => R1IN_4_3F(23),
  P(7) => R1IN_4_3F(24),
  P(8) => R1IN_4_3F(25),
  P(9) => R1IN_4_3F(26),
  P(10) => R1IN_4_3F(27),
  P(11) => R1IN_4_3F(28),
  P(12) => R1IN_4_3F(29),
  P(13) => R1IN_4_3F(30),
  P(14) => R1IN_4_3F(31),
  P(15) => R1IN_4_3F(32),
  P(16) => R1IN_4_3F(33),
  P(17) => R1IN_4_3F(34),
  P(18) => R1IN_4_3F(35),
  P(19) => R1IN_4_3F(36),
  P(20) => R1IN_4_3F(37),
  P(21) => R1IN_4_3F(38),
  P(22) => R1IN_4_3F(39),
  P(23) => R1IN_4_3F(40),
  P(24) => R1IN_4_3F(41),
  P(25) => R1IN_4_3F(42),
  P(26) => R1IN_4_3F(43),
  P(27) => UC_82,
  P(28) => UC_83,
  P(29) => UC_84,
  P(30) => UC_85,
  P(31) => UC_86,
  P(32) => UC_87,
  P(33) => UC_88,
  P(34) => UC_89,
  P(35) => UC_90,
  P(36) => UC_91,
  P(37) => UC_92,
  P(38) => UC_93,
  P(39) => UC_94,
  P(40) => UC_95,
  P(41) => UC_96,
  P(42) => UC_97,
  P(43) => UC_98,
  P(44) => UC_99,
  P(45) => UC_100,
  P(46) => UC_101,
  P(47) => UC_102,
  PCOUT(0) => R1IN_4_3_ADD_1_PCOUT(0),
  PCOUT(1) => R1IN_4_3_ADD_1_PCOUT(1),
  PCOUT(2) => R1IN_4_3_ADD_1_PCOUT(2),
  PCOUT(3) => R1IN_4_3_ADD_1_PCOUT(3),
  PCOUT(4) => R1IN_4_3_ADD_1_PCOUT(4),
  PCOUT(5) => R1IN_4_3_ADD_1_PCOUT(5),
  PCOUT(6) => R1IN_4_3_ADD_1_PCOUT(6),
  PCOUT(7) => R1IN_4_3_ADD_1_PCOUT(7),
  PCOUT(8) => R1IN_4_3_ADD_1_PCOUT(8),
  PCOUT(9) => R1IN_4_3_ADD_1_PCOUT(9),
  PCOUT(10) => R1IN_4_3_ADD_1_PCOUT(10),
  PCOUT(11) => R1IN_4_3_ADD_1_PCOUT(11),
  PCOUT(12) => R1IN_4_3_ADD_1_PCOUT(12),
  PCOUT(13) => R1IN_4_3_ADD_1_PCOUT(13),
  PCOUT(14) => R1IN_4_3_ADD_1_PCOUT(14),
  PCOUT(15) => R1IN_4_3_ADD_1_PCOUT(15),
  PCOUT(16) => R1IN_4_3_ADD_1_PCOUT(16),
  PCOUT(17) => R1IN_4_3_ADD_1_PCOUT(17),
  PCOUT(18) => R1IN_4_3_ADD_1_PCOUT(18),
  PCOUT(19) => R1IN_4_3_ADD_1_PCOUT(19),
  PCOUT(20) => R1IN_4_3_ADD_1_PCOUT(20),
  PCOUT(21) => R1IN_4_3_ADD_1_PCOUT(21),
  PCOUT(22) => R1IN_4_3_ADD_1_PCOUT(22),
  PCOUT(23) => R1IN_4_3_ADD_1_PCOUT(23),
  PCOUT(24) => R1IN_4_3_ADD_1_PCOUT(24),
  PCOUT(25) => R1IN_4_3_ADD_1_PCOUT(25),
  PCOUT(26) => R1IN_4_3_ADD_1_PCOUT(26),
  PCOUT(27) => R1IN_4_3_ADD_1_PCOUT(27),
  PCOUT(28) => R1IN_4_3_ADD_1_PCOUT(28),
  PCOUT(29) => R1IN_4_3_ADD_1_PCOUT(29),
  PCOUT(30) => R1IN_4_3_ADD_1_PCOUT(30),
  PCOUT(31) => R1IN_4_3_ADD_1_PCOUT(31),
  PCOUT(32) => R1IN_4_3_ADD_1_PCOUT(32),
  PCOUT(33) => R1IN_4_3_ADD_1_PCOUT(33),
  PCOUT(34) => R1IN_4_3_ADD_1_PCOUT(34),
  PCOUT(35) => R1IN_4_3_ADD_1_PCOUT(35),
  PCOUT(36) => R1IN_4_3_ADD_1_PCOUT(36),
  PCOUT(37) => R1IN_4_3_ADD_1_PCOUT(37),
  PCOUT(38) => R1IN_4_3_ADD_1_PCOUT(38),
  PCOUT(39) => R1IN_4_3_ADD_1_PCOUT(39),
  PCOUT(40) => R1IN_4_3_ADD_1_PCOUT(40),
  PCOUT(41) => R1IN_4_3_ADD_1_PCOUT(41),
  PCOUT(42) => R1IN_4_3_ADD_1_PCOUT(42),
  PCOUT(43) => R1IN_4_3_ADD_1_PCOUT(43),
  PCOUT(44) => R1IN_4_3_ADD_1_PCOUT(44),
  PCOUT(45) => R1IN_4_3_ADD_1_PCOUT(45),
  PCOUT(46) => R1IN_4_3_ADD_1_PCOUT(46),
  PCOUT(47) => R1IN_4_3_ADD_1_PCOUT(47));
R1IN_4_2_ADD_1q260w: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 1,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => A(51),
  A(1) => A(52),
  A(2) => A(53),
  A(3) => A(54),
  A(4) => A(55),
  A(5) => A(56),
  A(6) => A(57),
  A(7) => A(58),
  A(8) => A(59),
  A(9) => A(60),
  A(10) => NN_1,
  A(11) => NN_1,
  A(12) => NN_1,
  A(13) => NN_1,
  A(14) => NN_1,
  A(15) => NN_1,
  A(16) => NN_1,
  A(17) => NN_1,
  B(0) => B(17),
  B(1) => B(18),
  B(2) => B(19),
  B(3) => B(20),
  B(4) => B(21),
  B(5) => B(22),
  B(6) => B(23),
  B(7) => B(24),
  B(8) => B(25),
  B(9) => B(26),
  B(10) => B(27),
  B(11) => B(28),
  B(12) => B(29),
  B(13) => B(30),
  B(14) => B(31),
  B(15) => B(32),
  B(16) => B(33),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => R1IN_4_2_0(0),
  PCIN(1) => R1IN_4_2_0(1),
  PCIN(2) => R1IN_4_2_0(2),
  PCIN(3) => R1IN_4_2_0(3),
  PCIN(4) => R1IN_4_2_0(4),
  PCIN(5) => R1IN_4_2_0(5),
  PCIN(6) => R1IN_4_2_0(6),
  PCIN(7) => R1IN_4_2_0(7),
  PCIN(8) => R1IN_4_2_0(8),
  PCIN(9) => R1IN_4_2_0(9),
  PCIN(10) => R1IN_4_2_0(10),
  PCIN(11) => R1IN_4_2_0(11),
  PCIN(12) => R1IN_4_2_0(12),
  PCIN(13) => R1IN_4_2_0(13),
  PCIN(14) => R1IN_4_2_0(14),
  PCIN(15) => R1IN_4_2_0(15),
  PCIN(16) => R1IN_4_2_0(16),
  PCIN(17) => R1IN_4_2_1_0(17),
  PCIN(18) => R1IN_4_2_1_0(18),
  PCIN(19) => R1IN_4_2_1_0(19),
  PCIN(20) => R1IN_4_2_1_0(20),
  PCIN(21) => R1IN_4_2_1_0(21),
  PCIN(22) => R1IN_4_2_1_0(22),
  PCIN(23) => R1IN_4_2_1_0(23),
  PCIN(24) => R1IN_4_2_1_0(24),
  PCIN(25) => R1IN_4_2_1_0(25),
  PCIN(26) => R1IN_4_2_1_0(26),
  PCIN(27) => R1IN_4_2_1_0(27),
  PCIN(28) => R1IN_4_2_1_0(28),
  PCIN(29) => R1IN_4_2_1_0(29),
  PCIN(30) => R1IN_4_2_1_0(30),
  PCIN(31) => R1IN_4_2_1_0(31),
  PCIN(32) => R1IN_4_2_1_0(32),
  PCIN(33) => R1IN_4_2_1_0(33),
  PCIN(34) => UC_152_0,
  PCIN(35) => UC_153_0,
  PCIN(36) => UC_154_0,
  PCIN(37) => UC_155_0,
  PCIN(38) => UC_156_0,
  PCIN(39) => UC_157_0,
  PCIN(40) => UC_158_0,
  PCIN(41) => UC_159_0,
  PCIN(42) => UC_160_0,
  PCIN(43) => UC_161_0,
  PCIN(44) => UC_162_0,
  PCIN(45) => UC_163_0,
  PCIN(46) => UC_164_0,
  PCIN(47) => UC_165_0,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_2,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_2,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => CLK,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => EN,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_4_2_ADD_1_BCOUT(0),
  BCOUT(1) => R1IN_4_2_ADD_1_BCOUT(1),
  BCOUT(2) => R1IN_4_2_ADD_1_BCOUT(2),
  BCOUT(3) => R1IN_4_2_ADD_1_BCOUT(3),
  BCOUT(4) => R1IN_4_2_ADD_1_BCOUT(4),
  BCOUT(5) => R1IN_4_2_ADD_1_BCOUT(5),
  BCOUT(6) => R1IN_4_2_ADD_1_BCOUT(6),
  BCOUT(7) => R1IN_4_2_ADD_1_BCOUT(7),
  BCOUT(8) => R1IN_4_2_ADD_1_BCOUT(8),
  BCOUT(9) => R1IN_4_2_ADD_1_BCOUT(9),
  BCOUT(10) => R1IN_4_2_ADD_1_BCOUT(10),
  BCOUT(11) => R1IN_4_2_ADD_1_BCOUT(11),
  BCOUT(12) => R1IN_4_2_ADD_1_BCOUT(12),
  BCOUT(13) => R1IN_4_2_ADD_1_BCOUT(13),
  BCOUT(14) => R1IN_4_2_ADD_1_BCOUT(14),
  BCOUT(15) => R1IN_4_2_ADD_1_BCOUT(15),
  BCOUT(16) => R1IN_4_2_ADD_1_BCOUT(16),
  BCOUT(17) => R1IN_4_2_ADD_1_BCOUT(17),
  P(0) => R1IN_4_2F(17),
  P(1) => R1IN_4_2F(18),
  P(2) => R1IN_4_2F(19),
  P(3) => R1IN_4_2F(20),
  P(4) => R1IN_4_2F(21),
  P(5) => R1IN_4_2F(22),
  P(6) => R1IN_4_2F(23),
  P(7) => R1IN_4_2F(24),
  P(8) => R1IN_4_2F(25),
  P(9) => R1IN_4_2F(26),
  P(10) => R1IN_4_2F(27),
  P(11) => R1IN_4_2F(28),
  P(12) => R1IN_4_2F(29),
  P(13) => R1IN_4_2F(30),
  P(14) => R1IN_4_2F(31),
  P(15) => R1IN_4_2F(32),
  P(16) => R1IN_4_2F(33),
  P(17) => R1IN_4_2F(34),
  P(18) => R1IN_4_2F(35),
  P(19) => R1IN_4_2F(36),
  P(20) => R1IN_4_2F(37),
  P(21) => R1IN_4_2F(38),
  P(22) => R1IN_4_2F(39),
  P(23) => R1IN_4_2F(40),
  P(24) => R1IN_4_2F(41),
  P(25) => R1IN_4_2F(42),
  P(26) => R1IN_4_2F(43),
  P(27) => UC_61,
  P(28) => UC_62,
  P(29) => UC_63,
  P(30) => UC_64,
  P(31) => UC_65,
  P(32) => UC_66,
  P(33) => UC_67,
  P(34) => UC_68,
  P(35) => UC_69,
  P(36) => UC_70,
  P(37) => UC_71,
  P(38) => UC_72,
  P(39) => UC_73,
  P(40) => UC_74,
  P(41) => UC_75,
  P(42) => UC_76,
  P(43) => UC_77,
  P(44) => UC_78,
  P(45) => UC_79,
  P(46) => UC_80,
  P(47) => UC_81,
  PCOUT(0) => R1IN_4_2_ADD_1_PCOUT(0),
  PCOUT(1) => R1IN_4_2_ADD_1_PCOUT(1),
  PCOUT(2) => R1IN_4_2_ADD_1_PCOUT(2),
  PCOUT(3) => R1IN_4_2_ADD_1_PCOUT(3),
  PCOUT(4) => R1IN_4_2_ADD_1_PCOUT(4),
  PCOUT(5) => R1IN_4_2_ADD_1_PCOUT(5),
  PCOUT(6) => R1IN_4_2_ADD_1_PCOUT(6),
  PCOUT(7) => R1IN_4_2_ADD_1_PCOUT(7),
  PCOUT(8) => R1IN_4_2_ADD_1_PCOUT(8),
  PCOUT(9) => R1IN_4_2_ADD_1_PCOUT(9),
  PCOUT(10) => R1IN_4_2_ADD_1_PCOUT(10),
  PCOUT(11) => R1IN_4_2_ADD_1_PCOUT(11),
  PCOUT(12) => R1IN_4_2_ADD_1_PCOUT(12),
  PCOUT(13) => R1IN_4_2_ADD_1_PCOUT(13),
  PCOUT(14) => R1IN_4_2_ADD_1_PCOUT(14),
  PCOUT(15) => R1IN_4_2_ADD_1_PCOUT(15),
  PCOUT(16) => R1IN_4_2_ADD_1_PCOUT(16),
  PCOUT(17) => R1IN_4_2_ADD_1_PCOUT(17),
  PCOUT(18) => R1IN_4_2_ADD_1_PCOUT(18),
  PCOUT(19) => R1IN_4_2_ADD_1_PCOUT(19),
  PCOUT(20) => R1IN_4_2_ADD_1_PCOUT(20),
  PCOUT(21) => R1IN_4_2_ADD_1_PCOUT(21),
  PCOUT(22) => R1IN_4_2_ADD_1_PCOUT(22),
  PCOUT(23) => R1IN_4_2_ADD_1_PCOUT(23),
  PCOUT(24) => R1IN_4_2_ADD_1_PCOUT(24),
  PCOUT(25) => R1IN_4_2_ADD_1_PCOUT(25),
  PCOUT(26) => R1IN_4_2_ADD_1_PCOUT(26),
  PCOUT(27) => R1IN_4_2_ADD_1_PCOUT(27),
  PCOUT(28) => R1IN_4_2_ADD_1_PCOUT(28),
  PCOUT(29) => R1IN_4_2_ADD_1_PCOUT(29),
  PCOUT(30) => R1IN_4_2_ADD_1_PCOUT(30),
  PCOUT(31) => R1IN_4_2_ADD_1_PCOUT(31),
  PCOUT(32) => R1IN_4_2_ADD_1_PCOUT(32),
  PCOUT(33) => R1IN_4_2_ADD_1_PCOUT(33),
  PCOUT(34) => R1IN_4_2_ADD_1_PCOUT(34),
  PCOUT(35) => R1IN_4_2_ADD_1_PCOUT(35),
  PCOUT(36) => R1IN_4_2_ADD_1_PCOUT(36),
  PCOUT(37) => R1IN_4_2_ADD_1_PCOUT(37),
  PCOUT(38) => R1IN_4_2_ADD_1_PCOUT(38),
  PCOUT(39) => R1IN_4_2_ADD_1_PCOUT(39),
  PCOUT(40) => R1IN_4_2_ADD_1_PCOUT(40),
  PCOUT(41) => R1IN_4_2_ADD_1_PCOUT(41),
  PCOUT(42) => R1IN_4_2_ADD_1_PCOUT(42),
  PCOUT(43) => R1IN_4_2_ADD_1_PCOUT(43),
  PCOUT(44) => R1IN_4_2_ADD_1_PCOUT(44),
  PCOUT(45) => R1IN_4_2_ADD_1_PCOUT(45),
  PCOUT(46) => R1IN_4_2_ADD_1_PCOUT(46),
  PCOUT(47) => R1IN_4_2_ADD_1_PCOUT(47));
R1IN_3_2_ADD_1q260w: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 1,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => B(51),
  A(1) => B(52),
  A(2) => B(53),
  A(3) => B(54),
  A(4) => B(55),
  A(5) => B(56),
  A(6) => B(57),
  A(7) => B(58),
  A(8) => B(59),
  A(9) => B(60),
  A(10) => NN_1,
  A(11) => NN_1,
  A(12) => NN_1,
  A(13) => NN_1,
  A(14) => NN_1,
  A(15) => NN_1,
  A(16) => NN_1,
  A(17) => NN_1,
  B(0) => A(0),
  B(1) => A(1),
  B(2) => A(2),
  B(3) => A(3),
  B(4) => A(4),
  B(5) => A(5),
  B(6) => A(6),
  B(7) => A(7),
  B(8) => A(8),
  B(9) => A(9),
  B(10) => A(10),
  B(11) => A(11),
  B(12) => A(12),
  B(13) => A(13),
  B(14) => A(14),
  B(15) => A(15),
  B(16) => A(16),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => R1IN_3_2_0(0),
  PCIN(1) => R1IN_3_2_0(1),
  PCIN(2) => R1IN_3_2_0(2),
  PCIN(3) => R1IN_3_2_0(3),
  PCIN(4) => R1IN_3_2_0(4),
  PCIN(5) => R1IN_3_2_0(5),
  PCIN(6) => R1IN_3_2_0(6),
  PCIN(7) => R1IN_3_2_0(7),
  PCIN(8) => R1IN_3_2_0(8),
  PCIN(9) => R1IN_3_2_0(9),
  PCIN(10) => R1IN_3_2_0(10),
  PCIN(11) => R1IN_3_2_0(11),
  PCIN(12) => R1IN_3_2_0(12),
  PCIN(13) => R1IN_3_2_0(13),
  PCIN(14) => R1IN_3_2_0(14),
  PCIN(15) => R1IN_3_2_0(15),
  PCIN(16) => R1IN_3_2_0(16),
  PCIN(17) => R1IN_3_2_1_0(17),
  PCIN(18) => R1IN_3_2_1_0(18),
  PCIN(19) => R1IN_3_2_1_0(19),
  PCIN(20) => R1IN_3_2_1_0(20),
  PCIN(21) => R1IN_3_2_1_0(21),
  PCIN(22) => R1IN_3_2_1_0(22),
  PCIN(23) => R1IN_3_2_1_0(23),
  PCIN(24) => R1IN_3_2_1_0(24),
  PCIN(25) => R1IN_3_2_1_0(25),
  PCIN(26) => R1IN_3_2_1_0(26),
  PCIN(27) => R1IN_3_2_1_0(27),
  PCIN(28) => R1IN_3_2_1_0(28),
  PCIN(29) => R1IN_3_2_1_0(29),
  PCIN(30) => R1IN_3_2_1_0(30),
  PCIN(31) => R1IN_3_2_1_0(31),
  PCIN(32) => R1IN_3_2_1_0(32),
  PCIN(33) => R1IN_3_2_1_0(33),
  PCIN(34) => UC_138_0,
  PCIN(35) => UC_139_0,
  PCIN(36) => UC_140_0,
  PCIN(37) => UC_141_0,
  PCIN(38) => UC_142_0,
  PCIN(39) => UC_143_0,
  PCIN(40) => UC_144_0,
  PCIN(41) => UC_145_0,
  PCIN(42) => UC_146_0,
  PCIN(43) => UC_147_0,
  PCIN(44) => UC_148_0,
  PCIN(45) => UC_149_0,
  PCIN(46) => UC_150_0,
  PCIN(47) => UC_151_0,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_2,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_2,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => CLK,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => EN,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_3_2_ADD_1_BCOUT(0),
  BCOUT(1) => R1IN_3_2_ADD_1_BCOUT(1),
  BCOUT(2) => R1IN_3_2_ADD_1_BCOUT(2),
  BCOUT(3) => R1IN_3_2_ADD_1_BCOUT(3),
  BCOUT(4) => R1IN_3_2_ADD_1_BCOUT(4),
  BCOUT(5) => R1IN_3_2_ADD_1_BCOUT(5),
  BCOUT(6) => R1IN_3_2_ADD_1_BCOUT(6),
  BCOUT(7) => R1IN_3_2_ADD_1_BCOUT(7),
  BCOUT(8) => R1IN_3_2_ADD_1_BCOUT(8),
  BCOUT(9) => R1IN_3_2_ADD_1_BCOUT(9),
  BCOUT(10) => R1IN_3_2_ADD_1_BCOUT(10),
  BCOUT(11) => R1IN_3_2_ADD_1_BCOUT(11),
  BCOUT(12) => R1IN_3_2_ADD_1_BCOUT(12),
  BCOUT(13) => R1IN_3_2_ADD_1_BCOUT(13),
  BCOUT(14) => R1IN_3_2_ADD_1_BCOUT(14),
  BCOUT(15) => R1IN_3_2_ADD_1_BCOUT(15),
  BCOUT(16) => R1IN_3_2_ADD_1_BCOUT(16),
  BCOUT(17) => R1IN_3_2_ADD_1_BCOUT(17),
  P(0) => R1IN_3_2F(17),
  P(1) => R1IN_3_2F(18),
  P(2) => R1IN_3_2F(19),
  P(3) => R1IN_3_2F(20),
  P(4) => R1IN_3_2F(21),
  P(5) => R1IN_3_2F(22),
  P(6) => R1IN_3_2F(23),
  P(7) => R1IN_3_2F(24),
  P(8) => R1IN_3_2F(25),
  P(9) => R1IN_3_2F(26),
  P(10) => R1IN_3_2F(27),
  P(11) => R1IN_3_2F(28),
  P(12) => R1IN_3_2F(29),
  P(13) => R1IN_3_2F(30),
  P(14) => R1IN_3_2F(31),
  P(15) => R1IN_3_2F(32),
  P(16) => R1IN_3_2F(33),
  P(17) => R1IN_3_2F(34),
  P(18) => R1IN_3_2F(35),
  P(19) => R1IN_3_2F(36),
  P(20) => R1IN_3_2F(37),
  P(21) => R1IN_3_2F(38),
  P(22) => R1IN_3_2F(39),
  P(23) => R1IN_3_2F(40),
  P(24) => R1IN_3_2F(41),
  P(25) => R1IN_3_2F(42),
  P(26) => R1IN_3_2F(43),
  P(27) => UC_40,
  P(28) => UC_41,
  P(29) => UC_42,
  P(30) => UC_43,
  P(31) => UC_44,
  P(32) => UC_45,
  P(33) => UC_46,
  P(34) => UC_47,
  P(35) => UC_48,
  P(36) => UC_49,
  P(37) => UC_50,
  P(38) => UC_51,
  P(39) => UC_52,
  P(40) => UC_53,
  P(41) => UC_54,
  P(42) => UC_55,
  P(43) => UC_56,
  P(44) => UC_57,
  P(45) => UC_58,
  P(46) => UC_59,
  P(47) => UC_60,
  PCOUT(0) => R1IN_3_2_ADD_1_PCOUT(0),
  PCOUT(1) => R1IN_3_2_ADD_1_PCOUT(1),
  PCOUT(2) => R1IN_3_2_ADD_1_PCOUT(2),
  PCOUT(3) => R1IN_3_2_ADD_1_PCOUT(3),
  PCOUT(4) => R1IN_3_2_ADD_1_PCOUT(4),
  PCOUT(5) => R1IN_3_2_ADD_1_PCOUT(5),
  PCOUT(6) => R1IN_3_2_ADD_1_PCOUT(6),
  PCOUT(7) => R1IN_3_2_ADD_1_PCOUT(7),
  PCOUT(8) => R1IN_3_2_ADD_1_PCOUT(8),
  PCOUT(9) => R1IN_3_2_ADD_1_PCOUT(9),
  PCOUT(10) => R1IN_3_2_ADD_1_PCOUT(10),
  PCOUT(11) => R1IN_3_2_ADD_1_PCOUT(11),
  PCOUT(12) => R1IN_3_2_ADD_1_PCOUT(12),
  PCOUT(13) => R1IN_3_2_ADD_1_PCOUT(13),
  PCOUT(14) => R1IN_3_2_ADD_1_PCOUT(14),
  PCOUT(15) => R1IN_3_2_ADD_1_PCOUT(15),
  PCOUT(16) => R1IN_3_2_ADD_1_PCOUT(16),
  PCOUT(17) => R1IN_3_2_ADD_1_PCOUT(17),
  PCOUT(18) => R1IN_3_2_ADD_1_PCOUT(18),
  PCOUT(19) => R1IN_3_2_ADD_1_PCOUT(19),
  PCOUT(20) => R1IN_3_2_ADD_1_PCOUT(20),
  PCOUT(21) => R1IN_3_2_ADD_1_PCOUT(21),
  PCOUT(22) => R1IN_3_2_ADD_1_PCOUT(22),
  PCOUT(23) => R1IN_3_2_ADD_1_PCOUT(23),
  PCOUT(24) => R1IN_3_2_ADD_1_PCOUT(24),
  PCOUT(25) => R1IN_3_2_ADD_1_PCOUT(25),
  PCOUT(26) => R1IN_3_2_ADD_1_PCOUT(26),
  PCOUT(27) => R1IN_3_2_ADD_1_PCOUT(27),
  PCOUT(28) => R1IN_3_2_ADD_1_PCOUT(28),
  PCOUT(29) => R1IN_3_2_ADD_1_PCOUT(29),
  PCOUT(30) => R1IN_3_2_ADD_1_PCOUT(30),
  PCOUT(31) => R1IN_3_2_ADD_1_PCOUT(31),
  PCOUT(32) => R1IN_3_2_ADD_1_PCOUT(32),
  PCOUT(33) => R1IN_3_2_ADD_1_PCOUT(33),
  PCOUT(34) => R1IN_3_2_ADD_1_PCOUT(34),
  PCOUT(35) => R1IN_3_2_ADD_1_PCOUT(35),
  PCOUT(36) => R1IN_3_2_ADD_1_PCOUT(36),
  PCOUT(37) => R1IN_3_2_ADD_1_PCOUT(37),
  PCOUT(38) => R1IN_3_2_ADD_1_PCOUT(38),
  PCOUT(39) => R1IN_3_2_ADD_1_PCOUT(39),
  PCOUT(40) => R1IN_3_2_ADD_1_PCOUT(40),
  PCOUT(41) => R1IN_3_2_ADD_1_PCOUT(41),
  PCOUT(42) => R1IN_3_2_ADD_1_PCOUT(42),
  PCOUT(43) => R1IN_3_2_ADD_1_PCOUT(43),
  PCOUT(44) => R1IN_3_2_ADD_1_PCOUT(44),
  PCOUT(45) => R1IN_3_2_ADD_1_PCOUT(45),
  PCOUT(46) => R1IN_3_2_ADD_1_PCOUT(46),
  PCOUT(47) => R1IN_3_2_ADD_1_PCOUT(47));
R1IN_2_2_ADD_1q260w: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 1,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => A(51),
  A(1) => A(52),
  A(2) => A(53),
  A(3) => A(54),
  A(4) => A(55),
  A(5) => A(56),
  A(6) => A(57),
  A(7) => A(58),
  A(8) => A(59),
  A(9) => A(60),
  A(10) => NN_1,
  A(11) => NN_1,
  A(12) => NN_1,
  A(13) => NN_1,
  A(14) => NN_1,
  A(15) => NN_1,
  A(16) => NN_1,
  A(17) => NN_1,
  B(0) => B(0),
  B(1) => B(1),
  B(2) => B(2),
  B(3) => B(3),
  B(4) => B(4),
  B(5) => B(5),
  B(6) => B(6),
  B(7) => B(7),
  B(8) => B(8),
  B(9) => B(9),
  B(10) => B(10),
  B(11) => B(11),
  B(12) => B(12),
  B(13) => B(13),
  B(14) => B(14),
  B(15) => B(15),
  B(16) => B(16),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => R1IN_2_2_0(0),
  PCIN(1) => R1IN_2_2_0(1),
  PCIN(2) => R1IN_2_2_0(2),
  PCIN(3) => R1IN_2_2_0(3),
  PCIN(4) => R1IN_2_2_0(4),
  PCIN(5) => R1IN_2_2_0(5),
  PCIN(6) => R1IN_2_2_0(6),
  PCIN(7) => R1IN_2_2_0(7),
  PCIN(8) => R1IN_2_2_0(8),
  PCIN(9) => R1IN_2_2_0(9),
  PCIN(10) => R1IN_2_2_0(10),
  PCIN(11) => R1IN_2_2_0(11),
  PCIN(12) => R1IN_2_2_0(12),
  PCIN(13) => R1IN_2_2_0(13),
  PCIN(14) => R1IN_2_2_0(14),
  PCIN(15) => R1IN_2_2_0(15),
  PCIN(16) => R1IN_2_2_0(16),
  PCIN(17) => R1IN_2_2_1_0(17),
  PCIN(18) => R1IN_2_2_1_0(18),
  PCIN(19) => R1IN_2_2_1_0(19),
  PCIN(20) => R1IN_2_2_1_0(20),
  PCIN(21) => R1IN_2_2_1_0(21),
  PCIN(22) => R1IN_2_2_1_0(22),
  PCIN(23) => R1IN_2_2_1_0(23),
  PCIN(24) => R1IN_2_2_1_0(24),
  PCIN(25) => R1IN_2_2_1_0(25),
  PCIN(26) => R1IN_2_2_1_0(26),
  PCIN(27) => R1IN_2_2_1_0(27),
  PCIN(28) => R1IN_2_2_1_0(28),
  PCIN(29) => R1IN_2_2_1_0(29),
  PCIN(30) => R1IN_2_2_1_0(30),
  PCIN(31) => R1IN_2_2_1_0(31),
  PCIN(32) => R1IN_2_2_1_0(32),
  PCIN(33) => R1IN_2_2_1_0(33),
  PCIN(34) => UC_124_0,
  PCIN(35) => UC_125_0,
  PCIN(36) => UC_126_0,
  PCIN(37) => UC_127_0,
  PCIN(38) => UC_128_0,
  PCIN(39) => UC_129_0,
  PCIN(40) => UC_130_0,
  PCIN(41) => UC_131_0,
  PCIN(42) => UC_132_0,
  PCIN(43) => UC_133_0,
  PCIN(44) => UC_134_0,
  PCIN(45) => UC_135_0,
  PCIN(46) => UC_136_0,
  PCIN(47) => UC_137_0,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_2,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_2,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => CLK,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => EN,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_2_2_ADD_1_BCOUT(0),
  BCOUT(1) => R1IN_2_2_ADD_1_BCOUT(1),
  BCOUT(2) => R1IN_2_2_ADD_1_BCOUT(2),
  BCOUT(3) => R1IN_2_2_ADD_1_BCOUT(3),
  BCOUT(4) => R1IN_2_2_ADD_1_BCOUT(4),
  BCOUT(5) => R1IN_2_2_ADD_1_BCOUT(5),
  BCOUT(6) => R1IN_2_2_ADD_1_BCOUT(6),
  BCOUT(7) => R1IN_2_2_ADD_1_BCOUT(7),
  BCOUT(8) => R1IN_2_2_ADD_1_BCOUT(8),
  BCOUT(9) => R1IN_2_2_ADD_1_BCOUT(9),
  BCOUT(10) => R1IN_2_2_ADD_1_BCOUT(10),
  BCOUT(11) => R1IN_2_2_ADD_1_BCOUT(11),
  BCOUT(12) => R1IN_2_2_ADD_1_BCOUT(12),
  BCOUT(13) => R1IN_2_2_ADD_1_BCOUT(13),
  BCOUT(14) => R1IN_2_2_ADD_1_BCOUT(14),
  BCOUT(15) => R1IN_2_2_ADD_1_BCOUT(15),
  BCOUT(16) => R1IN_2_2_ADD_1_BCOUT(16),
  BCOUT(17) => R1IN_2_2_ADD_1_BCOUT(17),
  P(0) => R1IN_2_2F(17),
  P(1) => R1IN_2_2F(18),
  P(2) => R1IN_2_2F(19),
  P(3) => R1IN_2_2F(20),
  P(4) => R1IN_2_2F(21),
  P(5) => R1IN_2_2F(22),
  P(6) => R1IN_2_2F(23),
  P(7) => R1IN_2_2F(24),
  P(8) => R1IN_2_2F(25),
  P(9) => R1IN_2_2F(26),
  P(10) => R1IN_2_2F(27),
  P(11) => R1IN_2_2F(28),
  P(12) => R1IN_2_2F(29),
  P(13) => R1IN_2_2F(30),
  P(14) => R1IN_2_2F(31),
  P(15) => R1IN_2_2F(32),
  P(16) => R1IN_2_2F(33),
  P(17) => R1IN_2_2F(34),
  P(18) => R1IN_2_2F(35),
  P(19) => R1IN_2_2F(36),
  P(20) => R1IN_2_2F(37),
  P(21) => R1IN_2_2F(38),
  P(22) => R1IN_2_2F(39),
  P(23) => R1IN_2_2F(40),
  P(24) => R1IN_2_2F(41),
  P(25) => R1IN_2_2F(42),
  P(26) => R1IN_2_2F(43),
  P(27) => UC_19,
  P(28) => UC_20,
  P(29) => UC_21,
  P(30) => UC_22,
  P(31) => UC_23,
  P(32) => UC_24,
  P(33) => UC_25,
  P(34) => UC_26,
  P(35) => UC_27,
  P(36) => UC_28,
  P(37) => UC_29,
  P(38) => UC_30,
  P(39) => UC_31,
  P(40) => UC_32,
  P(41) => UC_33,
  P(42) => UC_34,
  P(43) => UC_35,
  P(44) => UC_36,
  P(45) => UC_37,
  P(46) => UC_38,
  P(47) => UC_39,
  PCOUT(0) => R1IN_2_2_ADD_1_PCOUT(0),
  PCOUT(1) => R1IN_2_2_ADD_1_PCOUT(1),
  PCOUT(2) => R1IN_2_2_ADD_1_PCOUT(2),
  PCOUT(3) => R1IN_2_2_ADD_1_PCOUT(3),
  PCOUT(4) => R1IN_2_2_ADD_1_PCOUT(4),
  PCOUT(5) => R1IN_2_2_ADD_1_PCOUT(5),
  PCOUT(6) => R1IN_2_2_ADD_1_PCOUT(6),
  PCOUT(7) => R1IN_2_2_ADD_1_PCOUT(7),
  PCOUT(8) => R1IN_2_2_ADD_1_PCOUT(8),
  PCOUT(9) => R1IN_2_2_ADD_1_PCOUT(9),
  PCOUT(10) => R1IN_2_2_ADD_1_PCOUT(10),
  PCOUT(11) => R1IN_2_2_ADD_1_PCOUT(11),
  PCOUT(12) => R1IN_2_2_ADD_1_PCOUT(12),
  PCOUT(13) => R1IN_2_2_ADD_1_PCOUT(13),
  PCOUT(14) => R1IN_2_2_ADD_1_PCOUT(14),
  PCOUT(15) => R1IN_2_2_ADD_1_PCOUT(15),
  PCOUT(16) => R1IN_2_2_ADD_1_PCOUT(16),
  PCOUT(17) => R1IN_2_2_ADD_1_PCOUT(17),
  PCOUT(18) => R1IN_2_2_ADD_1_PCOUT(18),
  PCOUT(19) => R1IN_2_2_ADD_1_PCOUT(19),
  PCOUT(20) => R1IN_2_2_ADD_1_PCOUT(20),
  PCOUT(21) => R1IN_2_2_ADD_1_PCOUT(21),
  PCOUT(22) => R1IN_2_2_ADD_1_PCOUT(22),
  PCOUT(23) => R1IN_2_2_ADD_1_PCOUT(23),
  PCOUT(24) => R1IN_2_2_ADD_1_PCOUT(24),
  PCOUT(25) => R1IN_2_2_ADD_1_PCOUT(25),
  PCOUT(26) => R1IN_2_2_ADD_1_PCOUT(26),
  PCOUT(27) => R1IN_2_2_ADD_1_PCOUT(27),
  PCOUT(28) => R1IN_2_2_ADD_1_PCOUT(28),
  PCOUT(29) => R1IN_2_2_ADD_1_PCOUT(29),
  PCOUT(30) => R1IN_2_2_ADD_1_PCOUT(30),
  PCOUT(31) => R1IN_2_2_ADD_1_PCOUT(31),
  PCOUT(32) => R1IN_2_2_ADD_1_PCOUT(32),
  PCOUT(33) => R1IN_2_2_ADD_1_PCOUT(33),
  PCOUT(34) => R1IN_2_2_ADD_1_PCOUT(34),
  PCOUT(35) => R1IN_2_2_ADD_1_PCOUT(35),
  PCOUT(36) => R1IN_2_2_ADD_1_PCOUT(36),
  PCOUT(37) => R1IN_2_2_ADD_1_PCOUT(37),
  PCOUT(38) => R1IN_2_2_ADD_1_PCOUT(38),
  PCOUT(39) => R1IN_2_2_ADD_1_PCOUT(39),
  PCOUT(40) => R1IN_2_2_ADD_1_PCOUT(40),
  PCOUT(41) => R1IN_2_2_ADD_1_PCOUT(41),
  PCOUT(42) => R1IN_2_2_ADD_1_PCOUT(42),
  PCOUT(43) => R1IN_2_2_ADD_1_PCOUT(43),
  PCOUT(44) => R1IN_2_2_ADD_1_PCOUT(44),
  PCOUT(45) => R1IN_2_2_ADD_1_PCOUT(45),
  PCOUT(46) => R1IN_2_2_ADD_1_PCOUT(46),
  PCOUT(47) => R1IN_2_2_ADD_1_PCOUT(47));
R1IN_4_4_ADD_1q270w: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 1,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => B(51),
  A(1) => B(52),
  A(2) => B(53),
  A(3) => B(54),
  A(4) => B(55),
  A(5) => B(56),
  A(6) => B(57),
  A(7) => B(58),
  A(8) => B(59),
  A(9) => B(60),
  A(10) => NN_1,
  A(11) => NN_1,
  A(12) => NN_1,
  A(13) => NN_1,
  A(14) => NN_1,
  A(15) => NN_1,
  A(16) => NN_1,
  A(17) => NN_1,
  B(0) => A(34),
  B(1) => A(35),
  B(2) => A(36),
  B(3) => A(37),
  B(4) => A(38),
  B(5) => A(39),
  B(6) => A(40),
  B(7) => A(41),
  B(8) => A(42),
  B(9) => A(43),
  B(10) => A(44),
  B(11) => A(45),
  B(12) => A(46),
  B(13) => A(47),
  B(14) => A(48),
  B(15) => A(49),
  B(16) => A(50),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => R1IN_4_4_2_0(0),
  PCIN(1) => R1IN_4_4_2_0(1),
  PCIN(2) => R1IN_4_4_2_0(2),
  PCIN(3) => R1IN_4_4_2_0(3),
  PCIN(4) => R1IN_4_4_2_0(4),
  PCIN(5) => R1IN_4_4_2_0(5),
  PCIN(6) => R1IN_4_4_2_0(6),
  PCIN(7) => R1IN_4_4_2_0(7),
  PCIN(8) => R1IN_4_4_2_0(8),
  PCIN(9) => R1IN_4_4_2_0(9),
  PCIN(10) => R1IN_4_4_2_0(10),
  PCIN(11) => R1IN_4_4_2_0(11),
  PCIN(12) => R1IN_4_4_2_0(12),
  PCIN(13) => R1IN_4_4_2_0(13),
  PCIN(14) => R1IN_4_4_2_0(14),
  PCIN(15) => R1IN_4_4_2_0(15),
  PCIN(16) => R1IN_4_4_2_0(16),
  PCIN(17) => R1IN_4_4_2_0(17),
  PCIN(18) => R1IN_4_4_2_0(18),
  PCIN(19) => R1IN_4_4_2_0(19),
  PCIN(20) => R1IN_4_4_2_0(20),
  PCIN(21) => R1IN_4_4_2_0(21),
  PCIN(22) => R1IN_4_4_2_0(22),
  PCIN(23) => R1IN_4_4_2_0(23),
  PCIN(24) => R1IN_4_4_2_0(24),
  PCIN(25) => R1IN_4_4_2_0(25),
  PCIN(26) => R1IN_4_4_2_0(26),
  PCIN(27) => UC_103_0,
  PCIN(28) => UC_104_0,
  PCIN(29) => UC_105_0,
  PCIN(30) => UC_106_0,
  PCIN(31) => UC_107_0,
  PCIN(32) => UC_108_0,
  PCIN(33) => UC_109_0,
  PCIN(34) => UC_110_0,
  PCIN(35) => UC_111_0,
  PCIN(36) => UC_112_0,
  PCIN(37) => UC_113_0,
  PCIN(38) => UC_114_0,
  PCIN(39) => UC_115_0,
  PCIN(40) => UC_116_0,
  PCIN(41) => UC_117_0,
  PCIN(42) => UC_118_0,
  PCIN(43) => UC_119_0,
  PCIN(44) => UC_120_0,
  PCIN(45) => UC_121_0,
  PCIN(46) => UC_122_0,
  PCIN(47) => UC_123_0,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_2,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => CLK,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => EN,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_4_4_ADD_1_BCOUT(0),
  BCOUT(1) => R1IN_4_4_ADD_1_BCOUT(1),
  BCOUT(2) => R1IN_4_4_ADD_1_BCOUT(2),
  BCOUT(3) => R1IN_4_4_ADD_1_BCOUT(3),
  BCOUT(4) => R1IN_4_4_ADD_1_BCOUT(4),
  BCOUT(5) => R1IN_4_4_ADD_1_BCOUT(5),
  BCOUT(6) => R1IN_4_4_ADD_1_BCOUT(6),
  BCOUT(7) => R1IN_4_4_ADD_1_BCOUT(7),
  BCOUT(8) => R1IN_4_4_ADD_1_BCOUT(8),
  BCOUT(9) => R1IN_4_4_ADD_1_BCOUT(9),
  BCOUT(10) => R1IN_4_4_ADD_1_BCOUT(10),
  BCOUT(11) => R1IN_4_4_ADD_1_BCOUT(11),
  BCOUT(12) => R1IN_4_4_ADD_1_BCOUT(12),
  BCOUT(13) => R1IN_4_4_ADD_1_BCOUT(13),
  BCOUT(14) => R1IN_4_4_ADD_1_BCOUT(14),
  BCOUT(15) => R1IN_4_4_ADD_1_BCOUT(15),
  BCOUT(16) => R1IN_4_4_ADD_1_BCOUT(16),
  BCOUT(17) => R1IN_4_4_ADD_1_BCOUT(17),
  P(0) => R1IN_4_4_ADD_1F(0),
  P(1) => R1IN_4_4_ADD_1F(1),
  P(2) => R1IN_4_4_ADD_1F(2),
  P(3) => R1IN_4_4_ADD_1F(3),
  P(4) => R1IN_4_4_ADD_1F(4),
  P(5) => R1IN_4_4_ADD_1F(5),
  P(6) => R1IN_4_4_ADD_1F(6),
  P(7) => R1IN_4_4_ADD_1F(7),
  P(8) => R1IN_4_4_ADD_1F(8),
  P(9) => R1IN_4_4_ADD_1F(9),
  P(10) => R1IN_4_4_ADD_1F(10),
  P(11) => R1IN_4_4_ADD_1F(11),
  P(12) => R1IN_4_4_ADD_1F(12),
  P(13) => R1IN_4_4_ADD_1F(13),
  P(14) => R1IN_4_4_ADD_1F(14),
  P(15) => R1IN_4_4_ADD_1F(15),
  P(16) => R1IN_4_4_ADD_1F(16),
  P(17) => R1IN_4_4_ADD_1F(17),
  P(18) => R1IN_4_4_ADD_1F(18),
  P(19) => R1IN_4_4_ADD_1F(19),
  P(20) => R1IN_4_4_ADD_1F(20),
  P(21) => R1IN_4_4_ADD_1F(21),
  P(22) => R1IN_4_4_ADD_1F(22),
  P(23) => R1IN_4_4_ADD_1F(23),
  P(24) => R1IN_4_4_ADD_1F(24),
  P(25) => R1IN_4_4_ADD_1F(25),
  P(26) => R1IN_4_4_ADD_1F(26),
  P(27) => R1IN_4_4_ADD_1F(27),
  P(28) => UC,
  P(29) => UC_0,
  P(30) => UC_1,
  P(31) => UC_2,
  P(32) => UC_3,
  P(33) => UC_4,
  P(34) => UC_5,
  P(35) => UC_6,
  P(36) => UC_7,
  P(37) => UC_8,
  P(38) => UC_9,
  P(39) => UC_10,
  P(40) => UC_11,
  P(41) => UC_12,
  P(42) => UC_13,
  P(43) => UC_14,
  P(44) => UC_15,
  P(45) => UC_16,
  P(46) => UC_17,
  P(47) => UC_18,
  PCOUT(0) => R1IN_4_4_ADD_1_PCOUT(0),
  PCOUT(1) => R1IN_4_4_ADD_1_PCOUT(1),
  PCOUT(2) => R1IN_4_4_ADD_1_PCOUT(2),
  PCOUT(3) => R1IN_4_4_ADD_1_PCOUT(3),
  PCOUT(4) => R1IN_4_4_ADD_1_PCOUT(4),
  PCOUT(5) => R1IN_4_4_ADD_1_PCOUT(5),
  PCOUT(6) => R1IN_4_4_ADD_1_PCOUT(6),
  PCOUT(7) => R1IN_4_4_ADD_1_PCOUT(7),
  PCOUT(8) => R1IN_4_4_ADD_1_PCOUT(8),
  PCOUT(9) => R1IN_4_4_ADD_1_PCOUT(9),
  PCOUT(10) => R1IN_4_4_ADD_1_PCOUT(10),
  PCOUT(11) => R1IN_4_4_ADD_1_PCOUT(11),
  PCOUT(12) => R1IN_4_4_ADD_1_PCOUT(12),
  PCOUT(13) => R1IN_4_4_ADD_1_PCOUT(13),
  PCOUT(14) => R1IN_4_4_ADD_1_PCOUT(14),
  PCOUT(15) => R1IN_4_4_ADD_1_PCOUT(15),
  PCOUT(16) => R1IN_4_4_ADD_1_PCOUT(16),
  PCOUT(17) => R1IN_4_4_ADD_1_PCOUT(17),
  PCOUT(18) => R1IN_4_4_ADD_1_PCOUT(18),
  PCOUT(19) => R1IN_4_4_ADD_1_PCOUT(19),
  PCOUT(20) => R1IN_4_4_ADD_1_PCOUT(20),
  PCOUT(21) => R1IN_4_4_ADD_1_PCOUT(21),
  PCOUT(22) => R1IN_4_4_ADD_1_PCOUT(22),
  PCOUT(23) => R1IN_4_4_ADD_1_PCOUT(23),
  PCOUT(24) => R1IN_4_4_ADD_1_PCOUT(24),
  PCOUT(25) => R1IN_4_4_ADD_1_PCOUT(25),
  PCOUT(26) => R1IN_4_4_ADD_1_PCOUT(26),
  PCOUT(27) => R1IN_4_4_ADD_1_PCOUT(27),
  PCOUT(28) => R1IN_4_4_ADD_1_PCOUT(28),
  PCOUT(29) => R1IN_4_4_ADD_1_PCOUT(29),
  PCOUT(30) => R1IN_4_4_ADD_1_PCOUT(30),
  PCOUT(31) => R1IN_4_4_ADD_1_PCOUT(31),
  PCOUT(32) => R1IN_4_4_ADD_1_PCOUT(32),
  PCOUT(33) => R1IN_4_4_ADD_1_PCOUT(33),
  PCOUT(34) => R1IN_4_4_ADD_1_PCOUT(34),
  PCOUT(35) => R1IN_4_4_ADD_1_PCOUT(35),
  PCOUT(36) => R1IN_4_4_ADD_1_PCOUT(36),
  PCOUT(37) => R1IN_4_4_ADD_1_PCOUT(37),
  PCOUT(38) => R1IN_4_4_ADD_1_PCOUT(38),
  PCOUT(39) => R1IN_4_4_ADD_1_PCOUT(39),
  PCOUT(40) => R1IN_4_4_ADD_1_PCOUT(40),
  PCOUT(41) => R1IN_4_4_ADD_1_PCOUT(41),
  PCOUT(42) => R1IN_4_4_ADD_1_PCOUT(42),
  PCOUT(43) => R1IN_4_4_ADD_1_PCOUT(43),
  PCOUT(44) => R1IN_4_4_ADD_1_PCOUT(44),
  PCOUT(45) => R1IN_4_4_ADD_1_PCOUT(45),
  PCOUT(46) => R1IN_4_4_ADD_1_PCOUT(46),
  PCOUT(47) => R1IN_4_4_ADD_1_PCOUT(47));
II_GND: GND port map (
    G => NN_1);
II_VCC: VCC port map (
    P => NN_2);
PRODUCT(17) <= NN_3;
end beh;


library ieee;
use ieee.std_logic_1164.all;
library UNISIM;
use UNISIM.VCOMPONENTS.all;

entity virtex6_mul_61x61 is
port(
  A : in std_logic_vector(60 downto 0);
  B : in std_logic_vector(60 downto 0);
  EN :  in std_logic;
  CLK :  in std_logic;
  PRODUCT : out std_logic_vector(121 downto 0));
end virtex6_mul_61x61;

architecture beh of virtex6_mul_61x61 is
  signal R1IN_3_2_1 : std_logic_vector(33 downto 17);
  signal R1IN_3_2 : std_logic_vector(16 downto 0);
  signal R1IN_2_2_1 : std_logic_vector(33 downto 17);
  signal R1IN_2_2 : std_logic_vector(16 downto 0);
  signal R1IN_4_4_2 : std_logic_vector(26 downto 0);
  signal R1IN_3 : std_logic_vector(60 downto 17);
  signal R1IN_2 : std_logic_vector(60 downto 17);
  signal R1IN_ADD_1 : std_logic_vector(32 downto 0);
  signal R1IN_4_4 : std_logic_vector(53 downto 17);
  signal R1IN_4 : std_logic_vector(54 downto 17);
  signal R1IN_4_3_1 : std_logic_vector(33 downto 17);
  signal R1IN_4_3 : std_logic_vector(16 downto 0);
  signal R1IN_4_ADD_1 : std_logic_vector(35 downto 1);
  signal R1IN_4_2 : std_logic_vector(16 downto 0);
  signal R1IN_4_2_1 : std_logic_vector(33 downto 17);
  signal R1IN_4F : std_logic_vector(52 downto 0);
  signal R1IN_4_1F : std_logic_vector(33 downto 17);
  signal R1IN_4_4F : std_logic_vector(16 downto 0);
  signal R1IN_4_2F : std_logic_vector(43 downto 1);
  signal R1IN_4_3F : std_logic_vector(43 downto 0);
  signal R1IN_1FF : std_logic_vector(33 downto 18);
  signal R1IN_4FF : std_logic_vector(16 downto 0);
  signal R1IN_ADD_1FF : std_logic_vector(32 downto 0);
  signal R1IN_4_4_1F : std_logic_vector(33 downto 18);
  signal R1IN_4_4_4F : std_logic_vector(19 downto 0);
  signal R1IN_4_4_ADD_1F : std_logic_vector(27 downto 0);
  signal R1IN_2F : std_logic_vector(16 downto 0);
  signal R1IN_3F : std_logic_vector(16 downto 0);
  signal R1IN_2_2F : std_logic_vector(43 downto 1);
  signal R1IN_2_1F : std_logic_vector(33 downto 17);
  signal R1IN_3_2F : std_logic_vector(43 downto 1);
  signal R1IN_3_1F : std_logic_vector(33 downto 17);
  signal R1IN_4_4_ADD_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_4_4_ADD_1_PCOUT : std_logic_vector(47 downto 0);
  signal R1IN_2_2_ADD_1_PCOUT : std_logic_vector(47 downto 0);
  signal R1IN_3_2_ADD_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_3_2_ADD_1_PCOUT : std_logic_vector(47 downto 0);
  signal R1IN_4_2_ADD_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_4_2_ADD_1_PCOUT : std_logic_vector(47 downto 0);
  signal R1IN_4_3_ADD_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_4_3_ADD_1_PCOUT : std_logic_vector(47 downto 0);
  signal R1IN_2_2_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_3_2_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_4_2_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_4_3_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_1_PCOUT : std_logic_vector(47 downto 0);
  signal R1IN_2_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_2_1_PCOUT : std_logic_vector(47 downto 0);
  signal R1IN_3_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_3_1_PCOUT : std_logic_vector(47 downto 0);
  signal R1IN_4_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_4_1_PCOUT : std_logic_vector(47 downto 0);
  signal R1IN_4_4_1_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_4_4_1_PCOUT : std_logic_vector(47 downto 0);
  signal R1IN_4_4_2_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_4_4_4_BCOUT : std_logic_vector(17 downto 0);
  signal R1IN_4_4_4_PCOUT : std_logic_vector(47 downto 0);
  signal R1IN_2_2_0 : std_logic_vector(16 downto 0);
  signal R1IN_2_2_1_0 : std_logic_vector(33 downto 17);
  signal R1IN_3_2_0 : std_logic_vector(16 downto 0);
  signal R1IN_3_2_1_0 : std_logic_vector(33 downto 17);
  signal R1IN_4_2_0 : std_logic_vector(16 downto 0);
  signal R1IN_4_2_1_0 : std_logic_vector(33 downto 17);
  signal R1IN_4_3_0 : std_logic_vector(16 downto 0);
  signal R1IN_4_3_1_0 : std_logic_vector(33 downto 17);
  signal R1IN_4_4_2_0 : std_logic_vector(26 downto 0);
  signal B_0 : std_logic_vector(16 downto 0);
  signal R1IN_3F_0 : std_logic_vector(16 downto 0);
  signal R1IN_3_1F_0 : std_logic_vector(33 downto 17);
  signal R1IN_2F_0 : std_logic_vector(16 downto 0);
  signal R1IN_2_1F_0 : std_logic_vector(33 downto 17);
  signal NN_1 : std_logic ;
  signal NN_2 : std_logic ;
  signal NN_12 : std_logic ;
  signal R1IN_ADD_2_0 : std_logic ;
  signal R1IN_4_4_ADD_2 : std_logic ;
  signal R1IN_2_ADD_1 : std_logic ;
  signal R1IN_3_ADD_1 : std_logic ;
  signal UC : std_logic ;
  signal UC_0 : std_logic ;
  signal UC_1 : std_logic ;
  signal UC_2 : std_logic ;
  signal UC_3 : std_logic ;
  signal UC_4 : std_logic ;
  signal UC_5 : std_logic ;
  signal UC_6 : std_logic ;
  signal UC_7 : std_logic ;
  signal UC_8 : std_logic ;
  signal UC_9 : std_logic ;
  signal UC_10 : std_logic ;
  signal UC_11 : std_logic ;
  signal UC_12 : std_logic ;
  signal UC_13 : std_logic ;
  signal UC_14 : std_logic ;
  signal UC_15 : std_logic ;
  signal UC_16 : std_logic ;
  signal UC_17 : std_logic ;
  signal UC_18 : std_logic ;
  signal UC_19 : std_logic ;
  signal UC_20 : std_logic ;
  signal UC_21 : std_logic ;
  signal UC_22 : std_logic ;
  signal UC_23 : std_logic ;
  signal UC_24 : std_logic ;
  signal UC_25 : std_logic ;
  signal UC_26 : std_logic ;
  signal UC_27 : std_logic ;
  signal UC_28 : std_logic ;
  signal UC_29 : std_logic ;
  signal UC_30 : std_logic ;
  signal UC_31 : std_logic ;
  signal UC_32 : std_logic ;
  signal UC_33 : std_logic ;
  signal UC_34 : std_logic ;
  signal UC_35 : std_logic ;
  signal UC_36 : std_logic ;
  signal UC_37 : std_logic ;
  signal UC_38 : std_logic ;
  signal UC_39 : std_logic ;
  signal UC_40 : std_logic ;
  signal UC_41 : std_logic ;
  signal UC_42 : std_logic ;
  signal UC_43 : std_logic ;
  signal UC_44 : std_logic ;
  signal UC_45 : std_logic ;
  signal UC_46 : std_logic ;
  signal UC_47 : std_logic ;
  signal UC_48 : std_logic ;
  signal UC_49 : std_logic ;
  signal UC_50 : std_logic ;
  signal UC_51 : std_logic ;
  signal UC_52 : std_logic ;
  signal UC_53 : std_logic ;
  signal UC_54 : std_logic ;
  signal UC_55 : std_logic ;
  signal UC_56 : std_logic ;
  signal UC_57 : std_logic ;
  signal UC_58 : std_logic ;
  signal UC_59 : std_logic ;
  signal UC_60 : std_logic ;
  signal UC_61 : std_logic ;
  signal UC_62 : std_logic ;
  signal UC_63 : std_logic ;
  signal UC_64 : std_logic ;
  signal UC_65 : std_logic ;
  signal UC_66 : std_logic ;
  signal UC_67 : std_logic ;
  signal UC_68 : std_logic ;
  signal UC_69 : std_logic ;
  signal UC_70 : std_logic ;
  signal UC_71 : std_logic ;
  signal UC_72 : std_logic ;
  signal UC_73 : std_logic ;
  signal UC_74 : std_logic ;
  signal UC_75 : std_logic ;
  signal UC_76 : std_logic ;
  signal UC_77 : std_logic ;
  signal UC_78 : std_logic ;
  signal UC_79 : std_logic ;
  signal UC_80 : std_logic ;
  signal UC_81 : std_logic ;
  signal UC_82 : std_logic ;
  signal UC_83 : std_logic ;
  signal UC_84 : std_logic ;
  signal UC_85 : std_logic ;
  signal UC_86 : std_logic ;
  signal UC_87 : std_logic ;
  signal UC_88 : std_logic ;
  signal UC_89 : std_logic ;
  signal UC_90 : std_logic ;
  signal UC_91 : std_logic ;
  signal UC_92 : std_logic ;
  signal UC_93 : std_logic ;
  signal UC_94 : std_logic ;
  signal UC_95 : std_logic ;
  signal UC_96 : std_logic ;
  signal UC_97 : std_logic ;
  signal UC_98 : std_logic ;
  signal UC_99 : std_logic ;
  signal UC_100 : std_logic ;
  signal UC_101 : std_logic ;
  signal UC_102 : std_logic ;
  signal UC_103 : std_logic ;
  signal UC_104 : std_logic ;
  signal UC_105 : std_logic ;
  signal UC_106 : std_logic ;
  signal UC_107 : std_logic ;
  signal UC_108 : std_logic ;
  signal UC_109 : std_logic ;
  signal UC_110 : std_logic ;
  signal UC_111 : std_logic ;
  signal UC_112 : std_logic ;
  signal UC_113 : std_logic ;
  signal UC_114 : std_logic ;
  signal UC_115 : std_logic ;
  signal UC_116 : std_logic ;
  signal UC_117 : std_logic ;
  signal UC_118 : std_logic ;
  signal UC_119 : std_logic ;
  signal UC_120 : std_logic ;
  signal UC_121 : std_logic ;
  signal UC_122 : std_logic ;
  signal UC_123 : std_logic ;
  signal UC_124 : std_logic ;
  signal UC_125 : std_logic ;
  signal UC_126 : std_logic ;
  signal UC_127 : std_logic ;
  signal UC_128 : std_logic ;
  signal UC_129 : std_logic ;
  signal UC_130 : std_logic ;
  signal UC_131 : std_logic ;
  signal UC_132 : std_logic ;
  signal UC_133 : std_logic ;
  signal UC_134 : std_logic ;
  signal UC_135 : std_logic ;
  signal UC_136 : std_logic ;
  signal UC_137 : std_logic ;
  signal UC_138 : std_logic ;
  signal UC_139 : std_logic ;
  signal UC_140 : std_logic ;
  signal UC_141 : std_logic ;
  signal UC_142 : std_logic ;
  signal UC_143 : std_logic ;
  signal UC_144 : std_logic ;
  signal UC_145 : std_logic ;
  signal UC_146 : std_logic ;
  signal UC_147 : std_logic ;
  signal UC_148 : std_logic ;
  signal UC_149 : std_logic ;
  signal UC_150 : std_logic ;
  signal UC_151 : std_logic ;
  signal UC_152 : std_logic ;
  signal UC_153 : std_logic ;
  signal UC_154 : std_logic ;
  signal UC_155 : std_logic ;
  signal UC_156 : std_logic ;
  signal UC_157 : std_logic ;
  signal UC_158 : std_logic ;
  signal UC_159 : std_logic ;
  signal UC_160 : std_logic ;
  signal UC_161 : std_logic ;
  signal UC_162 : std_logic ;
  signal UC_163 : std_logic ;
  signal UC_164 : std_logic ;
  signal UC_165 : std_logic ;
  signal UC_166 : std_logic ;
  signal UC_167 : std_logic ;
  signal UC_168 : std_logic ;
  signal UC_169 : std_logic ;
  signal UC_170 : std_logic ;
  signal UC_171 : std_logic ;
  signal UC_172 : std_logic ;
  signal UC_201 : std_logic ;
  signal UC_202 : std_logic ;
  signal UC_203 : std_logic ;
  signal UC_204 : std_logic ;
  signal UC_205 : std_logic ;
  signal UC_206 : std_logic ;
  signal UC_207 : std_logic ;
  signal UC_208 : std_logic ;
  signal UC_209 : std_logic ;
  signal UC_210 : std_logic ;
  signal UC_211 : std_logic ;
  signal UC_212 : std_logic ;
  signal UC_213 : std_logic ;
  signal UC_214 : std_logic ;
  signal UC_215 : std_logic ;
  signal UC_216 : std_logic ;
  signal UC_217 : std_logic ;
  signal UC_218 : std_logic ;
  signal UC_219 : std_logic ;
  signal UC_220 : std_logic ;
  signal UC_221 : std_logic ;
  signal UC_222 : std_logic ;
  signal UC_223 : std_logic ;
  signal UC_224 : std_logic ;
  signal UC_225 : std_logic ;
  signal UC_226 : std_logic ;
  signal UC_227 : std_logic ;
  signal UC_228 : std_logic ;
  signal UC_229 : std_logic ;
  signal UC_230 : std_logic ;
  signal UC_231 : std_logic ;
  signal UC_232 : std_logic ;
  signal UC_233 : std_logic ;
  signal UC_234 : std_logic ;
  signal UC_235 : std_logic ;
  signal UC_236 : std_logic ;
  signal UC_237 : std_logic ;
  signal UC_238 : std_logic ;
  signal UC_239 : std_logic ;
  signal UC_240 : std_logic ;
  signal UC_241 : std_logic ;
  signal UC_242 : std_logic ;
  signal UC_243 : std_logic ;
  signal UC_244 : std_logic ;
  signal UC_245 : std_logic ;
  signal UC_246 : std_logic ;
  signal UC_247 : std_logic ;
  signal UC_248 : std_logic ;
  signal UC_249 : std_logic ;
  signal UC_250 : std_logic ;
  signal UC_251 : std_logic ;
  signal UC_252 : std_logic ;
  signal UC_253 : std_logic ;
  signal UC_254 : std_logic ;
  signal UC_255 : std_logic ;
  signal UC_256 : std_logic ;
  signal UC_257 : std_logic ;
  signal UC_258 : std_logic ;
  signal UC_259 : std_logic ;
  signal UC_260 : std_logic ;
  signal UC_261 : std_logic ;
  signal UC_262 : std_logic ;
  signal UC_263 : std_logic ;
  signal UC_264 : std_logic ;
  signal UC_265 : std_logic ;
  signal UC_266 : std_logic ;
  signal UC_267 : std_logic ;
  signal UC_268 : std_logic ;
  signal UC_269 : std_logic ;
  signal UC_270 : std_logic ;
  signal UC_271 : std_logic ;
  signal UC_272 : std_logic ;
  signal UC_273 : std_logic ;
  signal UC_274 : std_logic ;
  signal UC_275 : std_logic ;
  signal UC_276 : std_logic ;
  signal UC_277 : std_logic ;
  signal UC_103_0 : std_logic ;
  signal UC_104_0 : std_logic ;
  signal UC_105_0 : std_logic ;
  signal UC_106_0 : std_logic ;
  signal UC_107_0 : std_logic ;
  signal UC_108_0 : std_logic ;
  signal UC_109_0 : std_logic ;
  signal UC_110_0 : std_logic ;
  signal UC_111_0 : std_logic ;
  signal UC_112_0 : std_logic ;
  signal UC_113_0 : std_logic ;
  signal UC_114_0 : std_logic ;
  signal UC_115_0 : std_logic ;
  signal UC_116_0 : std_logic ;
  signal UC_117_0 : std_logic ;
  signal UC_118_0 : std_logic ;
  signal UC_119_0 : std_logic ;
  signal UC_120_0 : std_logic ;
  signal UC_121_0 : std_logic ;
  signal UC_122_0 : std_logic ;
  signal UC_123_0 : std_logic ;
  signal UC_124_0 : std_logic ;
  signal UC_125_0 : std_logic ;
  signal UC_126_0 : std_logic ;
  signal UC_127_0 : std_logic ;
  signal UC_128_0 : std_logic ;
  signal UC_129_0 : std_logic ;
  signal UC_130_0 : std_logic ;
  signal UC_131_0 : std_logic ;
  signal UC_132_0 : std_logic ;
  signal UC_133_0 : std_logic ;
  signal UC_134_0 : std_logic ;
  signal UC_135_0 : std_logic ;
  signal UC_136_0 : std_logic ;
  signal UC_137_0 : std_logic ;
  signal UC_138_0 : std_logic ;
  signal UC_139_0 : std_logic ;
  signal UC_140_0 : std_logic ;
  signal UC_141_0 : std_logic ;
  signal UC_142_0 : std_logic ;
  signal UC_143_0 : std_logic ;
  signal UC_144_0 : std_logic ;
  signal UC_145_0 : std_logic ;
  signal UC_146_0 : std_logic ;
  signal UC_147_0 : std_logic ;
  signal UC_148_0 : std_logic ;
  signal UC_149_0 : std_logic ;
  signal UC_150_0 : std_logic ;
  signal UC_151_0 : std_logic ;
  signal UC_152_0 : std_logic ;
  signal UC_153_0 : std_logic ;
  signal UC_154_0 : std_logic ;
  signal UC_155_0 : std_logic ;
  signal UC_156_0 : std_logic ;
  signal UC_157_0 : std_logic ;
  signal UC_158_0 : std_logic ;
  signal UC_229_0 : std_logic ;
  signal UC_230_0 : std_logic ;
  signal UC_231_0 : std_logic ;
  signal UC_232_0 : std_logic ;
  signal UC_233_0 : std_logic ;
  signal UC_234_0 : std_logic ;
  signal UC_235_0 : std_logic ;
  signal UC_236_0 : std_logic ;
  signal UC_237_0 : std_logic ;
  signal UC_238_0 : std_logic ;
  signal UC_239_0 : std_logic ;
  signal UC_240_0 : std_logic ;
  signal UC_241_0 : std_logic ;
  signal UC_242_0 : std_logic ;
  signal UC_243_0 : std_logic ;
  signal UC_244_0 : std_logic ;
  signal UC_245_0 : std_logic ;
  signal UC_246_0 : std_logic ;
  signal UC_247_0 : std_logic ;
  signal UC_248_0 : std_logic ;
  signal UC_249_0 : std_logic ;
  signal GND_0 : std_logic ;
  signal R1IN_ADD_1_1_S_21 : std_logic ;
  signal R1IN_ADD_1_1_S_22 : std_logic ;
  signal R1IN_ADD_1_1_S_23 : std_logic ;
  signal R1IN_ADD_1_1_S_24 : std_logic ;
  signal R1IN_ADD_1_1_S_25 : std_logic ;
  signal R1IN_ADD_1_1_S_26 : std_logic ;
  signal R1IN_ADD_1_1_S_27 : std_logic ;
  signal R1IN_ADD_1_1_S_28 : std_logic ;
  signal R1IN_ADD_1_1_CRY_28 : std_logic ;
  signal R1IN_ADD_2_0_CRY_52 : std_logic ;
  signal R1IN_ADD_2_1_S_1 : std_logic ;
  signal R1IN_ADD_2_1_S_2 : std_logic ;
  signal R1IN_ADD_2_1_S_3 : std_logic ;
  signal R1IN_ADD_2_1_S_4 : std_logic ;
  signal R1IN_ADD_2_1_S_5 : std_logic ;
  signal R1IN_ADD_2_1_S_6 : std_logic ;
  signal R1IN_ADD_2_1_S_7 : std_logic ;
  signal R1IN_ADD_2_1_S_8 : std_logic ;
  signal R1IN_ADD_2_1_S_9 : std_logic ;
  signal R1IN_ADD_2_1_S_10 : std_logic ;
  signal R1IN_ADD_2_1_S_11 : std_logic ;
  signal R1IN_ADD_2_1_S_12 : std_logic ;
  signal R1IN_ADD_2_1_S_13 : std_logic ;
  signal R1IN_ADD_2_1_S_14 : std_logic ;
  signal R1IN_ADD_2_1_S_15 : std_logic ;
  signal R1IN_ADD_2_1_S_16 : std_logic ;
  signal R1IN_ADD_2_1_S_17 : std_logic ;
  signal R1IN_ADD_2_1_S_18 : std_logic ;
  signal R1IN_ADD_2_1_S_19 : std_logic ;
  signal R1IN_ADD_2_1_S_20 : std_logic ;
  signal R1IN_ADD_2_1_S_21 : std_logic ;
  signal R1IN_ADD_2_1_S_22 : std_logic ;
  signal R1IN_ADD_2_1_S_23 : std_logic ;
  signal R1IN_ADD_2_1_S_24 : std_logic ;
  signal R1IN_ADD_2_1_S_25 : std_logic ;
  signal R1IN_ADD_2_1_S_26 : std_logic ;
  signal R1IN_ADD_2_1_S_27 : std_logic ;
  signal R1IN_ADD_2_1_S_28 : std_logic ;
  signal R1IN_ADD_2_1_S_29 : std_logic ;
  signal R1IN_ADD_2_1_S_30 : std_logic ;
  signal R1IN_ADD_2_1_S_31 : std_logic ;
  signal R1IN_ADD_2_1_S_32 : std_logic ;
  signal R1IN_ADD_2_1_S_33 : std_logic ;
  signal R1IN_ADD_2_1_S_34 : std_logic ;
  signal R1IN_ADD_2_1_S_35 : std_logic ;
  signal R1IN_ADD_2_1_S_36 : std_logic ;
  signal R1IN_ADD_2_1_S_37 : std_logic ;
  signal R1IN_ADD_2_1_S_38 : std_logic ;
  signal R1IN_ADD_2_1_S_39 : std_logic ;
  signal R1IN_ADD_2_1_S_40 : std_logic ;
  signal R1IN_ADD_2_1_S_41 : std_logic ;
  signal R1IN_ADD_2_1_S_42 : std_logic ;
  signal R1IN_ADD_2_1_S_43 : std_logic ;
  signal R1IN_ADD_2_1_S_44 : std_logic ;
  signal R1IN_ADD_2_1_S_45 : std_logic ;
  signal R1IN_ADD_2_1_S_46 : std_logic ;
  signal R1IN_ADD_2_1_S_47 : std_logic ;
  signal R1IN_ADD_2_1_S_48 : std_logic ;
  signal R1IN_ADD_2_1_S_49 : std_logic ;
  signal R1IN_ADD_2_1_S_50 : std_logic ;
  signal R1IN_ADD_2_1_S_51 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_0 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_1 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_1 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_2 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_2 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_3 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_3 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_4 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_4 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_5 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_5 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_6 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_6 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_7 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_7 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_8 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_8 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_9 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_9 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_10 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_10 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_11 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_11 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_12 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_12 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_13 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_13 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_14 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_14 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_15 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_15 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_16 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_16 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_17 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_17 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_18 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_18 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_19 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_19 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_20 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_20 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_21 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_21 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_22 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_22 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_23 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_23 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_24 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_24 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_25 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_25 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_26 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_26 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_27 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_27 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_28 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_28 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_29 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_29 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_30 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_30 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_31 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_31 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_32 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_32 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_33 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_33 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_34 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_34 : std_logic ;
  signal R1IN_4_ADD_2_0_AXB_35 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_0 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_1 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_1 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_2 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_2 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_3 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_3 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_4 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_4 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_5 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_5 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_6 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_6 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_7 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_7 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_8 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_8 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_9 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_9 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_10 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_10 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_11 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_11 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_12 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_12 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_13 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_13 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_14 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_14 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_15 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_15 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_16 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_16 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_17 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_17 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_18 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_18 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_19 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_19 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_20 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_20 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_21 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_21 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_22 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_22 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_23 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_23 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_24 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_24 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_25 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_25 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_26 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_26 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_27 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_27 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_28 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_28 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_29 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_29 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_30 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_30 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_31 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_31 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_32 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_32 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_33 : std_logic ;
  signal R1IN_4_ADD_2_1_CRY_33 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_34 : std_logic ;
  signal R1IN_ADD_2_0_CRY_0 : std_logic ;
  signal R1IN_ADD_2_0_AXB_1 : std_logic ;
  signal R1IN_ADD_2_0_CRY_1 : std_logic ;
  signal R1IN_ADD_2_0_AXB_2 : std_logic ;
  signal R1IN_ADD_2_0_CRY_2 : std_logic ;
  signal R1IN_ADD_2_0_AXB_3 : std_logic ;
  signal R1IN_ADD_2_0_CRY_3 : std_logic ;
  signal R1IN_ADD_2_0_AXB_4 : std_logic ;
  signal R1IN_ADD_2_0_CRY_4 : std_logic ;
  signal R1IN_ADD_2_0_AXB_5 : std_logic ;
  signal R1IN_ADD_2_0_CRY_5 : std_logic ;
  signal R1IN_ADD_2_0_AXB_6 : std_logic ;
  signal R1IN_ADD_2_0_CRY_6 : std_logic ;
  signal R1IN_ADD_2_0_AXB_7 : std_logic ;
  signal R1IN_ADD_2_0_CRY_7 : std_logic ;
  signal R1IN_ADD_2_0_AXB_8 : std_logic ;
  signal R1IN_ADD_2_0_CRY_8 : std_logic ;
  signal R1IN_ADD_2_0_AXB_9 : std_logic ;
  signal R1IN_ADD_2_0_CRY_9 : std_logic ;
  signal R1IN_ADD_2_0_AXB_10 : std_logic ;
  signal R1IN_ADD_2_0_CRY_10 : std_logic ;
  signal R1IN_ADD_2_0_AXB_11 : std_logic ;
  signal R1IN_ADD_2_0_CRY_11 : std_logic ;
  signal R1IN_ADD_2_0_AXB_12 : std_logic ;
  signal R1IN_ADD_2_0_CRY_12 : std_logic ;
  signal R1IN_ADD_2_0_AXB_13 : std_logic ;
  signal R1IN_ADD_2_0_CRY_13 : std_logic ;
  signal R1IN_ADD_2_0_AXB_14 : std_logic ;
  signal R1IN_ADD_2_0_CRY_14 : std_logic ;
  signal R1IN_ADD_2_0_AXB_15 : std_logic ;
  signal R1IN_ADD_2_0_CRY_15 : std_logic ;
  signal R1IN_ADD_2_0_AXB_16 : std_logic ;
  signal R1IN_ADD_2_0_CRY_16 : std_logic ;
  signal R1IN_ADD_2_0_AXB_17 : std_logic ;
  signal R1IN_ADD_2_0_CRY_17 : std_logic ;
  signal R1IN_ADD_2_0_AXB_18 : std_logic ;
  signal R1IN_ADD_2_0_CRY_18 : std_logic ;
  signal R1IN_ADD_2_0_AXB_19 : std_logic ;
  signal R1IN_ADD_2_0_CRY_19 : std_logic ;
  signal R1IN_ADD_2_0_AXB_20 : std_logic ;
  signal R1IN_ADD_2_0_CRY_20 : std_logic ;
  signal R1IN_ADD_2_0_AXB_21 : std_logic ;
  signal R1IN_ADD_2_0_CRY_21 : std_logic ;
  signal R1IN_ADD_2_0_AXB_22 : std_logic ;
  signal R1IN_ADD_2_0_CRY_22 : std_logic ;
  signal R1IN_ADD_2_0_AXB_23 : std_logic ;
  signal R1IN_ADD_2_0_CRY_23 : std_logic ;
  signal R1IN_ADD_2_0_AXB_24 : std_logic ;
  signal R1IN_ADD_2_0_CRY_24 : std_logic ;
  signal R1IN_ADD_2_0_AXB_25 : std_logic ;
  signal R1IN_ADD_2_0_CRY_25 : std_logic ;
  signal R1IN_ADD_2_0_AXB_26 : std_logic ;
  signal R1IN_ADD_2_0_CRY_26 : std_logic ;
  signal R1IN_ADD_2_0_AXB_27 : std_logic ;
  signal R1IN_ADD_2_0_CRY_27 : std_logic ;
  signal R1IN_ADD_2_0_AXB_28 : std_logic ;
  signal R1IN_ADD_2_0_CRY_28 : std_logic ;
  signal R1IN_ADD_2_0_AXB_29 : std_logic ;
  signal R1IN_ADD_2_0_CRY_29 : std_logic ;
  signal R1IN_ADD_2_0_AXB_30 : std_logic ;
  signal R1IN_ADD_2_0_CRY_30 : std_logic ;
  signal R1IN_ADD_2_0_AXB_31 : std_logic ;
  signal R1IN_ADD_2_0_CRY_31 : std_logic ;
  signal R1IN_ADD_2_0_AXB_32 : std_logic ;
  signal R1IN_ADD_2_0_CRY_32 : std_logic ;
  signal R1IN_ADD_2_0_AXB_33 : std_logic ;
  signal R1IN_ADD_2_0_CRY_33 : std_logic ;
  signal R1IN_ADD_2_0_AXB_34 : std_logic ;
  signal R1IN_ADD_2_0_CRY_34 : std_logic ;
  signal R1IN_ADD_2_0_AXB_35 : std_logic ;
  signal R1IN_ADD_2_0_CRY_35 : std_logic ;
  signal R1IN_ADD_2_0_AXB_36 : std_logic ;
  signal R1IN_ADD_2_0_CRY_36 : std_logic ;
  signal R1IN_ADD_2_0_AXB_37 : std_logic ;
  signal R1IN_ADD_2_0_CRY_37 : std_logic ;
  signal R1IN_ADD_2_0_AXB_38 : std_logic ;
  signal R1IN_ADD_2_0_CRY_38 : std_logic ;
  signal R1IN_ADD_2_0_AXB_39 : std_logic ;
  signal R1IN_ADD_2_0_CRY_39 : std_logic ;
  signal R1IN_ADD_2_0_AXB_40 : std_logic ;
  signal R1IN_ADD_2_0_CRY_40 : std_logic ;
  signal R1IN_ADD_2_0_AXB_41 : std_logic ;
  signal R1IN_ADD_2_0_CRY_41 : std_logic ;
  signal R1IN_ADD_2_0_AXB_42 : std_logic ;
  signal R1IN_ADD_2_0_CRY_42 : std_logic ;
  signal R1IN_ADD_2_0_AXB_43 : std_logic ;
  signal R1IN_ADD_2_0_CRY_43 : std_logic ;
  signal R1IN_ADD_2_0_AXB_44 : std_logic ;
  signal R1IN_ADD_2_0_CRY_44 : std_logic ;
  signal R1IN_ADD_2_0_AXB_45 : std_logic ;
  signal R1IN_ADD_2_0_CRY_45 : std_logic ;
  signal R1IN_ADD_2_0_AXB_46 : std_logic ;
  signal R1IN_ADD_2_0_CRY_46 : std_logic ;
  signal R1IN_ADD_2_0_AXB_47 : std_logic ;
  signal R1IN_ADD_2_0_CRY_47 : std_logic ;
  signal R1IN_ADD_2_0_AXB_48 : std_logic ;
  signal R1IN_ADD_2_0_CRY_48 : std_logic ;
  signal R1IN_ADD_2_0_AXB_49 : std_logic ;
  signal R1IN_ADD_2_0_CRY_49 : std_logic ;
  signal R1IN_ADD_2_0_AXB_50 : std_logic ;
  signal R1IN_ADD_2_0_CRY_50 : std_logic ;
  signal R1IN_ADD_2_0_AXB_51 : std_logic ;
  signal R1IN_ADD_2_0_CRY_51 : std_logic ;
  signal R1IN_ADD_2_0_AXB_52 : std_logic ;
  signal R1IN_ADD_2_1_AXB_0 : std_logic ;
  signal R1IN_ADD_2_1_CRY_0 : std_logic ;
  signal R1IN_ADD_2_1_AXB_1 : std_logic ;
  signal R1IN_ADD_2_1_CRY_1 : std_logic ;
  signal R1IN_ADD_2_1_AXB_2 : std_logic ;
  signal R1IN_ADD_2_1_CRY_2 : std_logic ;
  signal R1IN_ADD_2_1_AXB_3 : std_logic ;
  signal R1IN_ADD_2_1_CRY_3 : std_logic ;
  signal R1IN_ADD_2_1_AXB_4 : std_logic ;
  signal R1IN_ADD_2_1_CRY_4 : std_logic ;
  signal R1IN_ADD_2_1_AXB_5 : std_logic ;
  signal R1IN_ADD_2_1_CRY_5 : std_logic ;
  signal R1IN_ADD_2_1_AXB_6 : std_logic ;
  signal R1IN_ADD_2_1_CRY_6 : std_logic ;
  signal R1IN_ADD_2_1_AXB_7 : std_logic ;
  signal R1IN_ADD_2_1_CRY_7 : std_logic ;
  signal R1IN_ADD_2_1_AXB_8 : std_logic ;
  signal R1IN_ADD_2_1_CRY_8 : std_logic ;
  signal R1IN_ADD_2_1_AXB_9 : std_logic ;
  signal R1IN_ADD_2_1_CRY_9 : std_logic ;
  signal R1IN_ADD_2_1_AXB_10 : std_logic ;
  signal R1IN_ADD_2_1_CRY_10 : std_logic ;
  signal R1IN_ADD_2_1_AXB_11 : std_logic ;
  signal R1IN_ADD_2_1_CRY_11 : std_logic ;
  signal R1IN_ADD_2_1_AXB_12 : std_logic ;
  signal R1IN_ADD_2_1_CRY_12 : std_logic ;
  signal R1IN_ADD_2_1_AXB_13 : std_logic ;
  signal R1IN_ADD_2_1_CRY_13 : std_logic ;
  signal R1IN_ADD_2_1_AXB_14 : std_logic ;
  signal R1IN_ADD_2_1_CRY_14 : std_logic ;
  signal R1IN_ADD_2_1_AXB_15 : std_logic ;
  signal R1IN_ADD_2_1_CRY_15 : std_logic ;
  signal R1IN_ADD_2_1_AXB_16 : std_logic ;
  signal R1IN_ADD_2_1_CRY_16 : std_logic ;
  signal R1IN_ADD_2_1_AXB_17 : std_logic ;
  signal R1IN_ADD_2_1_CRY_17 : std_logic ;
  signal R1IN_ADD_2_1_AXB_18 : std_logic ;
  signal R1IN_ADD_2_1_CRY_18 : std_logic ;
  signal R1IN_ADD_2_1_AXB_19 : std_logic ;
  signal R1IN_ADD_2_1_CRY_19 : std_logic ;
  signal R1IN_ADD_2_1_AXB_20 : std_logic ;
  signal R1IN_ADD_2_1_CRY_20 : std_logic ;
  signal R1IN_ADD_2_1_AXB_21 : std_logic ;
  signal R1IN_ADD_2_1_CRY_21 : std_logic ;
  signal R1IN_ADD_2_1_AXB_22 : std_logic ;
  signal R1IN_ADD_2_1_CRY_22 : std_logic ;
  signal R1IN_ADD_2_1_AXB_23 : std_logic ;
  signal R1IN_ADD_2_1_CRY_23 : std_logic ;
  signal R1IN_ADD_2_1_AXB_24 : std_logic ;
  signal R1IN_ADD_2_1_CRY_24 : std_logic ;
  signal R1IN_ADD_2_1_AXB_25 : std_logic ;
  signal R1IN_ADD_2_1_CRY_25 : std_logic ;
  signal R1IN_ADD_2_1_AXB_26 : std_logic ;
  signal R1IN_ADD_2_1_CRY_26 : std_logic ;
  signal R1IN_ADD_2_1_AXB_27 : std_logic ;
  signal R1IN_ADD_2_1_CRY_27 : std_logic ;
  signal R1IN_ADD_2_1_AXB_28 : std_logic ;
  signal R1IN_ADD_2_1_CRY_28 : std_logic ;
  signal R1IN_ADD_2_1_AXB_29 : std_logic ;
  signal R1IN_ADD_2_1_CRY_29 : std_logic ;
  signal R1IN_ADD_2_1_AXB_30 : std_logic ;
  signal R1IN_ADD_2_1_CRY_30 : std_logic ;
  signal R1IN_ADD_2_1_AXB_31 : std_logic ;
  signal R1IN_ADD_2_1_CRY_31 : std_logic ;
  signal R1IN_ADD_2_1_AXB_32 : std_logic ;
  signal R1IN_ADD_2_1_CRY_32 : std_logic ;
  signal R1IN_ADD_2_1_AXB_33 : std_logic ;
  signal R1IN_ADD_2_1_CRY_33 : std_logic ;
  signal R1IN_ADD_2_1_AXB_34 : std_logic ;
  signal R1IN_ADD_2_1_CRY_34 : std_logic ;
  signal R1IN_ADD_2_1_AXB_35 : std_logic ;
  signal R1IN_ADD_2_1_CRY_35 : std_logic ;
  signal R1IN_ADD_2_1_AXB_36 : std_logic ;
  signal R1IN_ADD_2_1_CRY_36 : std_logic ;
  signal R1IN_ADD_2_1_AXB_37 : std_logic ;
  signal R1IN_ADD_2_1_CRY_37 : std_logic ;
  signal R1IN_ADD_2_1_AXB_38 : std_logic ;
  signal R1IN_ADD_2_1_CRY_38 : std_logic ;
  signal R1IN_ADD_2_1_AXB_39 : std_logic ;
  signal R1IN_ADD_2_1_CRY_39 : std_logic ;
  signal R1IN_ADD_2_1_AXB_40 : std_logic ;
  signal R1IN_ADD_2_1_CRY_40 : std_logic ;
  signal R1IN_ADD_2_1_AXB_41 : std_logic ;
  signal R1IN_ADD_2_1_CRY_41 : std_logic ;
  signal R1IN_ADD_2_1_AXB_42 : std_logic ;
  signal R1IN_ADD_2_1_CRY_42 : std_logic ;
  signal R1IN_ADD_2_1_AXB_43 : std_logic ;
  signal R1IN_ADD_2_1_CRY_43 : std_logic ;
  signal R1IN_ADD_2_1_AXB_44 : std_logic ;
  signal R1IN_ADD_2_1_CRY_44 : std_logic ;
  signal R1IN_ADD_2_1_AXB_45 : std_logic ;
  signal R1IN_ADD_2_1_CRY_45 : std_logic ;
  signal R1IN_ADD_2_1_AXB_46 : std_logic ;
  signal R1IN_ADD_2_1_CRY_46 : std_logic ;
  signal R1IN_ADD_2_1_AXB_47 : std_logic ;
  signal R1IN_ADD_2_1_CRY_47 : std_logic ;
  signal R1IN_ADD_2_1_AXB_48 : std_logic ;
  signal R1IN_ADD_2_1_CRY_48 : std_logic ;
  signal R1IN_ADD_2_1_AXB_49 : std_logic ;
  signal R1IN_ADD_2_1_CRY_49 : std_logic ;
  signal R1IN_ADD_2_1_AXB_50 : std_logic ;
  signal R1IN_ADD_2_1_CRY_50 : std_logic ;
  signal R1IN_ADD_2_1_AXB_51 : std_logic ;
  signal R1IN_ADD_2_1_0_S_1 : std_logic ;
  signal R1IN_ADD_2_1_0_S_2 : std_logic ;
  signal R1IN_ADD_2_1_0_S_3 : std_logic ;
  signal R1IN_ADD_2_1_0_S_4 : std_logic ;
  signal R1IN_ADD_2_1_0_S_5 : std_logic ;
  signal R1IN_ADD_2_1_0_S_6 : std_logic ;
  signal R1IN_ADD_2_1_0_S_7 : std_logic ;
  signal R1IN_ADD_2_1_0_S_8 : std_logic ;
  signal R1IN_ADD_2_1_0_S_9 : std_logic ;
  signal R1IN_ADD_2_1_0_S_10 : std_logic ;
  signal R1IN_ADD_2_1_0_S_11 : std_logic ;
  signal R1IN_ADD_2_1_0_S_12 : std_logic ;
  signal R1IN_ADD_2_1_0_S_13 : std_logic ;
  signal R1IN_ADD_2_1_0_S_14 : std_logic ;
  signal R1IN_ADD_2_1_0_S_15 : std_logic ;
  signal R1IN_ADD_2_1_0_S_16 : std_logic ;
  signal R1IN_ADD_2_1_0_S_17 : std_logic ;
  signal R1IN_ADD_2_1_0_S_18 : std_logic ;
  signal R1IN_ADD_2_1_0_S_19 : std_logic ;
  signal R1IN_ADD_2_1_0_S_20 : std_logic ;
  signal R1IN_ADD_2_1_0_S_21 : std_logic ;
  signal R1IN_ADD_2_1_0_S_22 : std_logic ;
  signal R1IN_ADD_2_1_0_S_23 : std_logic ;
  signal R1IN_ADD_2_1_0_S_24 : std_logic ;
  signal R1IN_ADD_2_1_0_S_25 : std_logic ;
  signal R1IN_ADD_2_1_0_S_26 : std_logic ;
  signal R1IN_ADD_2_1_0_S_27 : std_logic ;
  signal R1IN_ADD_2_1_0_S_28 : std_logic ;
  signal R1IN_ADD_2_1_0_S_29 : std_logic ;
  signal R1IN_ADD_2_1_0_S_30 : std_logic ;
  signal R1IN_ADD_2_1_0_S_31 : std_logic ;
  signal R1IN_ADD_2_1_0_S_32 : std_logic ;
  signal R1IN_ADD_2_1_0_S_33 : std_logic ;
  signal R1IN_ADD_2_1_0_S_34 : std_logic ;
  signal R1IN_ADD_2_1_0_S_35 : std_logic ;
  signal R1IN_ADD_2_1_0_S_36 : std_logic ;
  signal R1IN_ADD_2_1_0_S_37 : std_logic ;
  signal R1IN_ADD_2_1_0_S_38 : std_logic ;
  signal R1IN_ADD_2_1_0_S_39 : std_logic ;
  signal R1IN_ADD_2_1_0_S_40 : std_logic ;
  signal R1IN_ADD_2_1_0_S_41 : std_logic ;
  signal R1IN_ADD_2_1_0_S_42 : std_logic ;
  signal R1IN_ADD_2_1_0_S_43 : std_logic ;
  signal R1IN_ADD_2_1_0_S_44 : std_logic ;
  signal R1IN_ADD_2_1_0_S_45 : std_logic ;
  signal R1IN_ADD_2_1_0_S_46 : std_logic ;
  signal R1IN_ADD_2_1_0_S_47 : std_logic ;
  signal R1IN_ADD_2_1_0_S_48 : std_logic ;
  signal R1IN_ADD_2_1_0_S_49 : std_logic ;
  signal R1IN_ADD_2_1_0_S_50 : std_logic ;
  signal R1IN_ADD_2_1_0_S_51 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_0 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_0 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_1 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_1 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_2 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_2 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_3 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_3 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_4 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_4 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_5 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_5 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_6 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_6 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_7 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_7 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_8 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_8 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_9 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_9 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_10 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_10 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_11 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_11 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_12 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_12 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_13 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_13 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_14 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_14 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_15 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_15 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_16 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_16 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_17 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_17 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_18 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_18 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_19 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_19 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_20 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_20 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_21 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_21 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_22 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_22 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_23 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_23 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_24 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_24 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_25 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_25 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_26 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_26 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_27 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_27 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_28 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_28 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_29 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_29 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_30 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_30 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_31 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_31 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_32 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_32 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_33 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_33 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_34 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_34 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_35 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_35 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_36 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_36 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_37 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_37 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_38 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_38 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_39 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_39 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_40 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_40 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_41 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_41 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_42 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_42 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_43 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_43 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_44 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_44 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_45 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_45 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_46 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_46 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_47 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_47 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_48 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_48 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_49 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_49 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_50 : std_logic ;
  signal R1IN_ADD_2_1_0_CRY_50 : std_logic ;
  signal R1IN_ADD_2_1_0_AXB_51 : std_logic ;
  signal R1IN_ADD_1_0_CRY_0 : std_logic ;
  signal R1IN_ADD_1_0_AXB_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_1 : std_logic ;
  signal R1IN_ADD_1_0_AXB_2 : std_logic ;
  signal R1IN_ADD_1_0_CRY_2 : std_logic ;
  signal R1IN_ADD_1_0_AXB_3 : std_logic ;
  signal R1IN_ADD_1_0_CRY_3 : std_logic ;
  signal R1IN_ADD_1_0_AXB_4 : std_logic ;
  signal R1IN_ADD_1_0_CRY_4 : std_logic ;
  signal R1IN_ADD_1_0_AXB_5 : std_logic ;
  signal R1IN_ADD_1_0_CRY_5 : std_logic ;
  signal R1IN_ADD_1_0_AXB_6 : std_logic ;
  signal R1IN_ADD_1_0_CRY_6 : std_logic ;
  signal R1IN_ADD_1_0_AXB_7 : std_logic ;
  signal R1IN_ADD_1_0_CRY_7 : std_logic ;
  signal R1IN_ADD_1_0_AXB_8 : std_logic ;
  signal R1IN_ADD_1_0_CRY_8 : std_logic ;
  signal R1IN_ADD_1_0_AXB_9 : std_logic ;
  signal R1IN_ADD_1_0_CRY_9 : std_logic ;
  signal R1IN_ADD_1_0_AXB_10 : std_logic ;
  signal R1IN_ADD_1_0_CRY_10 : std_logic ;
  signal R1IN_ADD_1_0_AXB_11 : std_logic ;
  signal R1IN_ADD_1_0_CRY_11 : std_logic ;
  signal R1IN_ADD_1_0_AXB_12 : std_logic ;
  signal R1IN_ADD_1_0_CRY_12 : std_logic ;
  signal R1IN_ADD_1_0_AXB_13 : std_logic ;
  signal R1IN_ADD_1_0_CRY_13 : std_logic ;
  signal R1IN_ADD_1_0_AXB_14 : std_logic ;
  signal R1IN_ADD_1_0_CRY_14 : std_logic ;
  signal R1IN_ADD_1_0_AXB_15 : std_logic ;
  signal R1IN_ADD_1_0_CRY_15 : std_logic ;
  signal R1IN_ADD_1_0_AXB_16 : std_logic ;
  signal R1IN_ADD_1_0_CRY_16 : std_logic ;
  signal R1IN_ADD_1_0_AXB_17 : std_logic ;
  signal R1IN_ADD_1_0_CRY_17 : std_logic ;
  signal R1IN_ADD_1_0_AXB_18 : std_logic ;
  signal R1IN_ADD_1_0_CRY_18 : std_logic ;
  signal R1IN_ADD_1_0_AXB_19 : std_logic ;
  signal R1IN_ADD_1_0_CRY_19 : std_logic ;
  signal R1IN_ADD_1_0_AXB_20 : std_logic ;
  signal R1IN_ADD_1_0_CRY_20 : std_logic ;
  signal R1IN_ADD_1_0_AXB_21 : std_logic ;
  signal R1IN_ADD_1_0_CRY_21 : std_logic ;
  signal R1IN_ADD_1_0_AXB_22 : std_logic ;
  signal R1IN_ADD_1_0_CRY_22 : std_logic ;
  signal R1IN_ADD_1_0_AXB_23 : std_logic ;
  signal R1IN_ADD_1_0_CRY_23 : std_logic ;
  signal R1IN_ADD_1_0_AXB_24 : std_logic ;
  signal R1IN_ADD_1_0_CRY_24 : std_logic ;
  signal R1IN_ADD_1_0_AXB_25 : std_logic ;
  signal R1IN_ADD_1_0_CRY_25 : std_logic ;
  signal R1IN_ADD_1_0_AXB_26 : std_logic ;
  signal R1IN_ADD_1_0_CRY_26 : std_logic ;
  signal R1IN_ADD_1_0_AXB_27 : std_logic ;
  signal R1IN_ADD_1_0_CRY_27 : std_logic ;
  signal R1IN_ADD_1_0_AXB_28 : std_logic ;
  signal R1IN_ADD_1_0_CRY_28 : std_logic ;
  signal R1IN_ADD_1_0_AXB_29 : std_logic ;
  signal R1IN_ADD_1_0_CRY_29 : std_logic ;
  signal R1IN_ADD_1_0_AXB_30 : std_logic ;
  signal R1IN_ADD_1_0_CRY_30 : std_logic ;
  signal R1IN_ADD_1_0_AXB_31 : std_logic ;
  signal R1IN_ADD_1_1_AXB_0 : std_logic ;
  signal R1IN_ADD_1_1_CRY_0 : std_logic ;
  signal R1IN_ADD_1_1_AXB_1 : std_logic ;
  signal R1IN_ADD_1_1_CRY_1 : std_logic ;
  signal R1IN_ADD_1_1_AXB_2 : std_logic ;
  signal R1IN_ADD_1_1_CRY_2 : std_logic ;
  signal R1IN_ADD_1_1_AXB_3 : std_logic ;
  signal R1IN_ADD_1_1_CRY_3 : std_logic ;
  signal R1IN_ADD_1_1_AXB_4 : std_logic ;
  signal R1IN_ADD_1_1_CRY_4 : std_logic ;
  signal R1IN_ADD_1_1_AXB_5 : std_logic ;
  signal R1IN_ADD_1_1_CRY_5 : std_logic ;
  signal R1IN_ADD_1_1_AXB_6 : std_logic ;
  signal R1IN_ADD_1_1_CRY_6 : std_logic ;
  signal R1IN_ADD_1_1_AXB_7 : std_logic ;
  signal R1IN_ADD_1_1_CRY_7 : std_logic ;
  signal R1IN_ADD_1_1_AXB_8 : std_logic ;
  signal R1IN_ADD_1_1_CRY_8 : std_logic ;
  signal R1IN_ADD_1_1_AXB_9 : std_logic ;
  signal R1IN_ADD_1_1_CRY_9 : std_logic ;
  signal R1IN_ADD_1_1_AXB_10 : std_logic ;
  signal R1IN_ADD_1_1_CRY_10 : std_logic ;
  signal R1IN_ADD_1_1_AXB_11 : std_logic ;
  signal R1IN_ADD_1_1_CRY_11 : std_logic ;
  signal R1IN_ADD_1_1_AXB_12 : std_logic ;
  signal R1IN_ADD_1_1_CRY_12 : std_logic ;
  signal R1IN_ADD_1_1_AXB_13 : std_logic ;
  signal R1IN_ADD_1_1_CRY_13 : std_logic ;
  signal R1IN_ADD_1_1_AXB_14 : std_logic ;
  signal R1IN_ADD_1_1_CRY_14 : std_logic ;
  signal R1IN_ADD_1_1_AXB_15 : std_logic ;
  signal R1IN_ADD_1_1_CRY_15 : std_logic ;
  signal R1IN_ADD_1_1_AXB_16 : std_logic ;
  signal R1IN_ADD_1_1_CRY_16 : std_logic ;
  signal R1IN_ADD_1_1_AXB_17 : std_logic ;
  signal R1IN_ADD_1_1_CRY_17 : std_logic ;
  signal R1IN_ADD_1_1_AXB_18 : std_logic ;
  signal R1IN_ADD_1_1_CRY_18 : std_logic ;
  signal R1IN_ADD_1_1_AXB_19 : std_logic ;
  signal R1IN_ADD_1_1_CRY_19 : std_logic ;
  signal R1IN_ADD_1_1_AXB_20 : std_logic ;
  signal R1IN_ADD_1_1_CRY_20 : std_logic ;
  signal R1IN_ADD_1_1_AXB_21 : std_logic ;
  signal R1IN_ADD_1_1_CRY_21 : std_logic ;
  signal R1IN_ADD_1_1_AXB_22 : std_logic ;
  signal R1IN_ADD_1_1_CRY_22 : std_logic ;
  signal R1IN_ADD_1_1_AXB_23 : std_logic ;
  signal R1IN_ADD_1_1_CRY_23 : std_logic ;
  signal R1IN_ADD_1_1_AXB_24 : std_logic ;
  signal R1IN_ADD_1_1_CRY_24 : std_logic ;
  signal R1IN_ADD_1_1_AXB_25 : std_logic ;
  signal R1IN_ADD_1_1_CRY_25 : std_logic ;
  signal R1IN_ADD_1_1_AXB_26 : std_logic ;
  signal R1IN_ADD_1_1_CRY_26 : std_logic ;
  signal R1IN_ADD_1_1_AXB_27 : std_logic ;
  signal R1IN_ADD_1_1_CRY_27 : std_logic ;
  signal R1IN_ADD_1_1_AXB_28 : std_logic ;
  signal R1IN_ADD_1_1_0_S_21 : std_logic ;
  signal R1IN_ADD_1_1_0_S_22 : std_logic ;
  signal R1IN_ADD_1_1_0_S_23 : std_logic ;
  signal R1IN_ADD_1_1_0_S_24 : std_logic ;
  signal R1IN_ADD_1_1_0_S_25 : std_logic ;
  signal R1IN_ADD_1_1_0_S_26 : std_logic ;
  signal R1IN_ADD_1_1_0_S_27 : std_logic ;
  signal R1IN_ADD_1_1_0_S_28 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_28 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_0 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_0 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_1 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_1 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_2 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_2 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_3 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_3 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_4 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_4 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_5 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_5 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_6 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_6 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_7 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_7 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_8 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_8 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_9 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_9 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_10 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_10 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_11 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_11 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_12 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_12 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_13 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_13 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_14 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_14 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_15 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_15 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_16 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_16 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_17 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_17 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_18 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_18 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_19 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_19 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_20 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_20 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_21 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_21 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_22 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_22 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_23 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_23 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_24 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_24 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_25 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_25 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_26 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_26 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_27 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_27 : std_logic ;
  signal R1IN_ADD_1_1_0_AXB_28 : std_logic ;
  signal R1IN_3_ADD_1_CRY_0 : std_logic ;
  signal R1IN_3_ADD_1_AXB_1 : std_logic ;
  signal R1IN_3_ADD_1_CRY_1 : std_logic ;
  signal R1IN_3_ADD_1_AXB_2 : std_logic ;
  signal R1IN_3_ADD_1_CRY_2 : std_logic ;
  signal R1IN_3_ADD_1_AXB_3 : std_logic ;
  signal R1IN_3_ADD_1_CRY_3 : std_logic ;
  signal R1IN_3_ADD_1_AXB_4 : std_logic ;
  signal R1IN_3_ADD_1_CRY_4 : std_logic ;
  signal R1IN_3_ADD_1_AXB_5 : std_logic ;
  signal R1IN_3_ADD_1_CRY_5 : std_logic ;
  signal R1IN_3_ADD_1_AXB_6 : std_logic ;
  signal R1IN_3_ADD_1_CRY_6 : std_logic ;
  signal R1IN_3_ADD_1_AXB_7 : std_logic ;
  signal R1IN_3_ADD_1_CRY_7 : std_logic ;
  signal R1IN_3_ADD_1_AXB_8 : std_logic ;
  signal R1IN_3_ADD_1_CRY_8 : std_logic ;
  signal R1IN_3_ADD_1_AXB_9 : std_logic ;
  signal R1IN_3_ADD_1_CRY_9 : std_logic ;
  signal R1IN_3_ADD_1_AXB_10 : std_logic ;
  signal R1IN_3_ADD_1_CRY_10 : std_logic ;
  signal R1IN_3_ADD_1_AXB_11 : std_logic ;
  signal R1IN_3_ADD_1_CRY_11 : std_logic ;
  signal R1IN_3_ADD_1_AXB_12 : std_logic ;
  signal R1IN_3_ADD_1_CRY_12 : std_logic ;
  signal R1IN_3_ADD_1_AXB_13 : std_logic ;
  signal R1IN_3_ADD_1_CRY_13 : std_logic ;
  signal R1IN_3_ADD_1_AXB_14 : std_logic ;
  signal R1IN_3_ADD_1_CRY_14 : std_logic ;
  signal R1IN_3_ADD_1_AXB_15 : std_logic ;
  signal R1IN_3_ADD_1_CRY_15 : std_logic ;
  signal R1IN_3_ADD_1_AXB_16 : std_logic ;
  signal R1IN_3_ADD_1_CRY_16 : std_logic ;
  signal R1IN_3_ADD_1_AXB_17 : std_logic ;
  signal R1IN_3_ADD_1_CRY_17 : std_logic ;
  signal R1IN_3_ADD_1_AXB_18 : std_logic ;
  signal R1IN_3_ADD_1_CRY_18 : std_logic ;
  signal R1IN_3_ADD_1_AXB_19 : std_logic ;
  signal R1IN_3_ADD_1_CRY_19 : std_logic ;
  signal R1IN_3_ADD_1_AXB_20 : std_logic ;
  signal R1IN_3_ADD_1_CRY_20 : std_logic ;
  signal R1IN_3_ADD_1_AXB_21 : std_logic ;
  signal R1IN_3_ADD_1_CRY_21 : std_logic ;
  signal R1IN_3_ADD_1_AXB_22 : std_logic ;
  signal R1IN_3_ADD_1_CRY_22 : std_logic ;
  signal R1IN_3_ADD_1_AXB_23 : std_logic ;
  signal R1IN_3_ADD_1_CRY_23 : std_logic ;
  signal R1IN_3_ADD_1_AXB_24 : std_logic ;
  signal R1IN_3_ADD_1_CRY_24 : std_logic ;
  signal R1IN_3_ADD_1_AXB_25 : std_logic ;
  signal R1IN_3_ADD_1_CRY_25 : std_logic ;
  signal R1IN_3_ADD_1_AXB_26 : std_logic ;
  signal R1IN_3_ADD_1_CRY_26 : std_logic ;
  signal R1IN_3_ADD_1_AXB_27 : std_logic ;
  signal R1IN_3_ADD_1_CRY_27 : std_logic ;
  signal R1IN_3_ADD_1_AXB_28 : std_logic ;
  signal R1IN_3_ADD_1_CRY_28 : std_logic ;
  signal R1IN_3_ADD_1_AXB_29 : std_logic ;
  signal R1IN_3_ADD_1_CRY_29 : std_logic ;
  signal R1IN_3_ADD_1_AXB_30 : std_logic ;
  signal R1IN_3_ADD_1_CRY_30 : std_logic ;
  signal R1IN_3_ADD_1_AXB_31 : std_logic ;
  signal R1IN_3_ADD_1_CRY_31 : std_logic ;
  signal R1IN_3_ADD_1_AXB_32 : std_logic ;
  signal R1IN_3_ADD_1_CRY_32 : std_logic ;
  signal R1IN_3_ADD_1_AXB_33 : std_logic ;
  signal R1IN_3_ADD_1_CRY_33 : std_logic ;
  signal R1IN_3_ADD_1_AXB_34 : std_logic ;
  signal R1IN_3_ADD_1_CRY_34 : std_logic ;
  signal R1IN_3_ADD_1_AXB_35 : std_logic ;
  signal R1IN_3_ADD_1_CRY_35 : std_logic ;
  signal R1IN_3_ADD_1_AXB_36 : std_logic ;
  signal R1IN_3_ADD_1_CRY_36 : std_logic ;
  signal R1IN_3_ADD_1_AXB_37 : std_logic ;
  signal R1IN_3_ADD_1_CRY_37 : std_logic ;
  signal R1IN_3_ADD_1_AXB_38 : std_logic ;
  signal R1IN_3_ADD_1_CRY_38 : std_logic ;
  signal R1IN_3_ADD_1_AXB_39 : std_logic ;
  signal R1IN_3_ADD_1_CRY_39 : std_logic ;
  signal R1IN_3_ADD_1_AXB_40 : std_logic ;
  signal R1IN_3_ADD_1_CRY_40 : std_logic ;
  signal R1IN_3_ADD_1_AXB_41 : std_logic ;
  signal R1IN_3_ADD_1_CRY_41 : std_logic ;
  signal R1IN_3_ADD_1_AXB_42 : std_logic ;
  signal R1IN_3_ADD_1_CRY_42 : std_logic ;
  signal R1IN_3_ADD_1_AXB_43 : std_logic ;
  signal R1IN_2_ADD_1_CRY_0 : std_logic ;
  signal R1IN_2_ADD_1_AXB_1 : std_logic ;
  signal R1IN_2_ADD_1_CRY_1 : std_logic ;
  signal R1IN_2_ADD_1_AXB_2 : std_logic ;
  signal R1IN_2_ADD_1_CRY_2 : std_logic ;
  signal R1IN_2_ADD_1_AXB_3 : std_logic ;
  signal R1IN_2_ADD_1_CRY_3 : std_logic ;
  signal R1IN_2_ADD_1_AXB_4 : std_logic ;
  signal R1IN_2_ADD_1_CRY_4 : std_logic ;
  signal R1IN_2_ADD_1_AXB_5 : std_logic ;
  signal R1IN_2_ADD_1_CRY_5 : std_logic ;
  signal R1IN_2_ADD_1_AXB_6 : std_logic ;
  signal R1IN_2_ADD_1_CRY_6 : std_logic ;
  signal R1IN_2_ADD_1_AXB_7 : std_logic ;
  signal R1IN_2_ADD_1_CRY_7 : std_logic ;
  signal R1IN_2_ADD_1_AXB_8 : std_logic ;
  signal R1IN_2_ADD_1_CRY_8 : std_logic ;
  signal R1IN_2_ADD_1_AXB_9 : std_logic ;
  signal R1IN_2_ADD_1_CRY_9 : std_logic ;
  signal R1IN_2_ADD_1_AXB_10 : std_logic ;
  signal R1IN_2_ADD_1_CRY_10 : std_logic ;
  signal R1IN_2_ADD_1_AXB_11 : std_logic ;
  signal R1IN_2_ADD_1_CRY_11 : std_logic ;
  signal R1IN_2_ADD_1_AXB_12 : std_logic ;
  signal R1IN_2_ADD_1_CRY_12 : std_logic ;
  signal R1IN_2_ADD_1_AXB_13 : std_logic ;
  signal R1IN_2_ADD_1_CRY_13 : std_logic ;
  signal R1IN_2_ADD_1_AXB_14 : std_logic ;
  signal R1IN_2_ADD_1_CRY_14 : std_logic ;
  signal R1IN_2_ADD_1_AXB_15 : std_logic ;
  signal R1IN_2_ADD_1_CRY_15 : std_logic ;
  signal R1IN_2_ADD_1_AXB_16 : std_logic ;
  signal R1IN_2_ADD_1_CRY_16 : std_logic ;
  signal R1IN_2_ADD_1_AXB_17 : std_logic ;
  signal R1IN_2_ADD_1_CRY_17 : std_logic ;
  signal R1IN_2_ADD_1_AXB_18 : std_logic ;
  signal R1IN_2_ADD_1_CRY_18 : std_logic ;
  signal R1IN_2_ADD_1_AXB_19 : std_logic ;
  signal R1IN_2_ADD_1_CRY_19 : std_logic ;
  signal R1IN_2_ADD_1_AXB_20 : std_logic ;
  signal R1IN_2_ADD_1_CRY_20 : std_logic ;
  signal R1IN_2_ADD_1_AXB_21 : std_logic ;
  signal R1IN_2_ADD_1_CRY_21 : std_logic ;
  signal R1IN_2_ADD_1_AXB_22 : std_logic ;
  signal R1IN_2_ADD_1_CRY_22 : std_logic ;
  signal R1IN_2_ADD_1_AXB_23 : std_logic ;
  signal R1IN_2_ADD_1_CRY_23 : std_logic ;
  signal R1IN_2_ADD_1_AXB_24 : std_logic ;
  signal R1IN_2_ADD_1_CRY_24 : std_logic ;
  signal R1IN_2_ADD_1_AXB_25 : std_logic ;
  signal R1IN_2_ADD_1_CRY_25 : std_logic ;
  signal R1IN_2_ADD_1_AXB_26 : std_logic ;
  signal R1IN_2_ADD_1_CRY_26 : std_logic ;
  signal R1IN_2_ADD_1_AXB_27 : std_logic ;
  signal R1IN_2_ADD_1_CRY_27 : std_logic ;
  signal R1IN_2_ADD_1_AXB_28 : std_logic ;
  signal R1IN_2_ADD_1_CRY_28 : std_logic ;
  signal R1IN_2_ADD_1_AXB_29 : std_logic ;
  signal R1IN_2_ADD_1_CRY_29 : std_logic ;
  signal R1IN_2_ADD_1_AXB_30 : std_logic ;
  signal R1IN_2_ADD_1_CRY_30 : std_logic ;
  signal R1IN_2_ADD_1_AXB_31 : std_logic ;
  signal R1IN_2_ADD_1_CRY_31 : std_logic ;
  signal R1IN_2_ADD_1_AXB_32 : std_logic ;
  signal R1IN_2_ADD_1_CRY_32 : std_logic ;
  signal R1IN_2_ADD_1_AXB_33 : std_logic ;
  signal R1IN_2_ADD_1_CRY_33 : std_logic ;
  signal R1IN_2_ADD_1_AXB_34 : std_logic ;
  signal R1IN_2_ADD_1_CRY_34 : std_logic ;
  signal R1IN_2_ADD_1_AXB_35 : std_logic ;
  signal R1IN_2_ADD_1_CRY_35 : std_logic ;
  signal R1IN_2_ADD_1_AXB_36 : std_logic ;
  signal R1IN_2_ADD_1_CRY_36 : std_logic ;
  signal R1IN_2_ADD_1_AXB_37 : std_logic ;
  signal R1IN_2_ADD_1_CRY_37 : std_logic ;
  signal R1IN_2_ADD_1_AXB_38 : std_logic ;
  signal R1IN_2_ADD_1_CRY_38 : std_logic ;
  signal R1IN_2_ADD_1_AXB_39 : std_logic ;
  signal R1IN_2_ADD_1_CRY_39 : std_logic ;
  signal R1IN_2_ADD_1_AXB_40 : std_logic ;
  signal R1IN_2_ADD_1_CRY_40 : std_logic ;
  signal R1IN_2_ADD_1_AXB_41 : std_logic ;
  signal R1IN_2_ADD_1_CRY_41 : std_logic ;
  signal R1IN_2_ADD_1_AXB_42 : std_logic ;
  signal R1IN_2_ADD_1_CRY_42 : std_logic ;
  signal R1IN_2_ADD_1_AXB_43 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_0 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_1 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_1 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_2 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_2 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_3 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_3 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_4 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_4 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_5 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_5 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_6 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_6 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_7 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_7 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_8 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_8 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_9 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_9 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_10 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_10 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_11 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_11 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_12 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_12 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_13 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_13 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_14 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_14 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_15 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_15 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_16 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_16 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_17 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_17 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_18 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_18 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_19 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_19 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_20 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_20 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_21 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_21 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_22 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_22 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_23 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_23 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_24 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_24 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_25 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_25 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_26 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_26 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_27 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_27 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_28 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_28 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_29 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_29 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_30 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_30 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_31 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_31 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_32 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_32 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_33 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_33 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_34 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_34 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_35 : std_logic ;
  signal R1IN_4_4_ADD_2_CRY_35 : std_logic ;
  signal R1IN_4_4_ADD_2_AXB_36 : std_logic ;
  signal R1IN_4_ADD_2_0 : std_logic ;
  signal R1IN_4_ADD_1_CRY_0 : std_logic ;
  signal R1IN_4_ADD_1_AXB_1 : std_logic ;
  signal R1IN_4_ADD_1_CRY_1 : std_logic ;
  signal R1IN_4_ADD_1_AXB_2 : std_logic ;
  signal R1IN_4_ADD_1_CRY_2 : std_logic ;
  signal R1IN_4_ADD_1_AXB_3 : std_logic ;
  signal R1IN_4_ADD_1_CRY_3 : std_logic ;
  signal R1IN_4_ADD_1_AXB_4 : std_logic ;
  signal R1IN_4_ADD_1_CRY_4 : std_logic ;
  signal R1IN_4_ADD_1_AXB_5 : std_logic ;
  signal R1IN_4_ADD_1_CRY_5 : std_logic ;
  signal R1IN_4_ADD_1_AXB_6 : std_logic ;
  signal R1IN_4_ADD_1_CRY_6 : std_logic ;
  signal R1IN_4_ADD_1_AXB_7 : std_logic ;
  signal R1IN_4_ADD_1_CRY_7 : std_logic ;
  signal R1IN_4_ADD_1_AXB_8 : std_logic ;
  signal R1IN_4_ADD_1_CRY_8 : std_logic ;
  signal R1IN_4_ADD_1_AXB_9 : std_logic ;
  signal R1IN_4_ADD_1_CRY_9 : std_logic ;
  signal R1IN_4_ADD_1_AXB_10 : std_logic ;
  signal R1IN_4_ADD_1_CRY_10 : std_logic ;
  signal R1IN_4_ADD_1_AXB_11 : std_logic ;
  signal R1IN_4_ADD_1_CRY_11 : std_logic ;
  signal R1IN_4_ADD_1_AXB_12 : std_logic ;
  signal R1IN_4_ADD_1_CRY_12 : std_logic ;
  signal R1IN_4_ADD_1_AXB_13 : std_logic ;
  signal R1IN_4_ADD_1_CRY_13 : std_logic ;
  signal R1IN_4_ADD_1_AXB_14 : std_logic ;
  signal R1IN_4_ADD_1_CRY_14 : std_logic ;
  signal R1IN_4_ADD_1_AXB_15 : std_logic ;
  signal R1IN_4_ADD_1_CRY_15 : std_logic ;
  signal R1IN_4_ADD_1_AXB_16 : std_logic ;
  signal R1IN_4_ADD_1_CRY_16 : std_logic ;
  signal R1IN_4_ADD_1_AXB_17 : std_logic ;
  signal R1IN_4_ADD_1_CRY_17 : std_logic ;
  signal R1IN_4_ADD_1_AXB_18 : std_logic ;
  signal R1IN_4_ADD_1_CRY_18 : std_logic ;
  signal R1IN_4_ADD_1_AXB_19 : std_logic ;
  signal R1IN_4_ADD_1_CRY_19 : std_logic ;
  signal R1IN_4_ADD_1_AXB_20 : std_logic ;
  signal R1IN_4_ADD_1_CRY_20 : std_logic ;
  signal R1IN_4_ADD_1_AXB_21 : std_logic ;
  signal R1IN_4_ADD_1_CRY_21 : std_logic ;
  signal R1IN_4_ADD_1_AXB_22 : std_logic ;
  signal R1IN_4_ADD_1_CRY_22 : std_logic ;
  signal R1IN_4_ADD_1_AXB_23 : std_logic ;
  signal R1IN_4_ADD_1_CRY_23 : std_logic ;
  signal R1IN_4_ADD_1_AXB_24 : std_logic ;
  signal R1IN_4_ADD_1_CRY_24 : std_logic ;
  signal R1IN_4_ADD_1_AXB_25 : std_logic ;
  signal R1IN_4_ADD_1_CRY_25 : std_logic ;
  signal R1IN_4_ADD_1_AXB_26 : std_logic ;
  signal R1IN_4_ADD_1_CRY_26 : std_logic ;
  signal R1IN_4_ADD_1_AXB_27 : std_logic ;
  signal R1IN_4_ADD_1_CRY_27 : std_logic ;
  signal R1IN_4_ADD_1_AXB_28 : std_logic ;
  signal R1IN_4_ADD_1_CRY_28 : std_logic ;
  signal R1IN_4_ADD_1_AXB_29 : std_logic ;
  signal R1IN_4_ADD_1_CRY_29 : std_logic ;
  signal R1IN_4_ADD_1_AXB_30 : std_logic ;
  signal R1IN_4_ADD_1_CRY_30 : std_logic ;
  signal R1IN_4_ADD_1_AXB_31 : std_logic ;
  signal R1IN_4_ADD_1_CRY_31 : std_logic ;
  signal R1IN_4_ADD_1_AXB_32 : std_logic ;
  signal R1IN_4_ADD_1_CRY_32 : std_logic ;
  signal R1IN_4_ADD_1_AXB_33 : std_logic ;
  signal R1IN_4_ADD_1_CRY_33 : std_logic ;
  signal R1IN_4_ADD_1_AXB_34 : std_logic ;
  signal R1IN_4_ADD_1_CRY_34 : std_logic ;
  signal R1IN_4_ADD_1_AXB_35 : std_logic ;
  signal R1IN_4_ADD_1_CRY_35 : std_logic ;
  signal R1IN_4_ADD_1_AXB_36 : std_logic ;
  signal R1IN_4_ADD_1_CRY_36 : std_logic ;
  signal R1IN_4_ADD_1_AXB_37 : std_logic ;
  signal R1IN_4_ADD_1_CRY_37 : std_logic ;
  signal R1IN_4_ADD_1_AXB_38 : std_logic ;
  signal R1IN_4_ADD_1_CRY_38 : std_logic ;
  signal R1IN_4_ADD_1_AXB_39 : std_logic ;
  signal R1IN_4_ADD_1_CRY_39 : std_logic ;
  signal R1IN_4_ADD_1_AXB_40 : std_logic ;
  signal R1IN_4_ADD_1_CRY_40 : std_logic ;
  signal R1IN_4_ADD_1_AXB_41 : std_logic ;
  signal R1IN_4_ADD_1_CRY_41 : std_logic ;
  signal R1IN_4_ADD_1_AXB_42 : std_logic ;
  signal R1IN_4_ADD_1_CRY_42 : std_logic ;
  signal R1IN_4_ADD_1_AXB_43 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO : std_logic ;
  signal N_5444 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_0 : std_logic ;
  signal N_5445 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_1 : std_logic ;
  signal N_5446 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_2 : std_logic ;
  signal N_5447 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_3 : std_logic ;
  signal N_5448 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_4 : std_logic ;
  signal N_5449 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_5 : std_logic ;
  signal N_5450 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_6 : std_logic ;
  signal N_5451 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_7 : std_logic ;
  signal N_5452 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_8 : std_logic ;
  signal N_5453 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_9 : std_logic ;
  signal N_5454 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_10 : std_logic ;
  signal N_5455 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_11 : std_logic ;
  signal N_5456 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_12 : std_logic ;
  signal N_5457 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_13 : std_logic ;
  signal N_5458 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_14 : std_logic ;
  signal N_5459 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_15 : std_logic ;
  signal N_5460 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_16 : std_logic ;
  signal N_5461 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_17 : std_logic ;
  signal N_5462 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_18 : std_logic ;
  signal N_5463 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_19 : std_logic ;
  signal N_5464 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_20 : std_logic ;
  signal N_5465 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_21 : std_logic ;
  signal N_5466 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_22 : std_logic ;
  signal N_5467 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_23 : std_logic ;
  signal N_5468 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_24 : std_logic ;
  signal N_5469 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_25 : std_logic ;
  signal N_5470 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_26 : std_logic ;
  signal N_5471 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_27 : std_logic ;
  signal N_5472 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_28 : std_logic ;
  signal N_5473 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_29 : std_logic ;
  signal N_5474 : std_logic ;
  signal N_1577 : std_logic ;
  signal R2_PIPE_157_RET : std_logic ;
  signal N_1913 : std_logic ;
  signal R2_PIPE_157_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO : std_logic ;
  signal N_5475 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_30 : std_logic ;
  signal N_5476 : std_logic ;
  signal N_1575 : std_logic ;
  signal R2_PIPE_156_RET : std_logic ;
  signal N_1912 : std_logic ;
  signal R2_PIPE_156_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_0 : std_logic ;
  signal N_5477 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_31 : std_logic ;
  signal N_5478 : std_logic ;
  signal N_1573 : std_logic ;
  signal R2_PIPE_155_RET : std_logic ;
  signal N_1911 : std_logic ;
  signal R2_PIPE_155_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_1 : std_logic ;
  signal N_5479 : std_logic ;
  signal N_1571 : std_logic ;
  signal R2_PIPE_154_RET : std_logic ;
  signal N_1910 : std_logic ;
  signal R2_PIPE_154_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_2 : std_logic ;
  signal N_5480 : std_logic ;
  signal N_1569 : std_logic ;
  signal R2_PIPE_153_RET : std_logic ;
  signal N_1909 : std_logic ;
  signal R2_PIPE_153_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_3 : std_logic ;
  signal N_5481 : std_logic ;
  signal N_1567 : std_logic ;
  signal R2_PIPE_152_RET : std_logic ;
  signal N_1908 : std_logic ;
  signal R2_PIPE_152_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_4 : std_logic ;
  signal N_5482 : std_logic ;
  signal N_1565 : std_logic ;
  signal R2_PIPE_151_RET : std_logic ;
  signal N_1907 : std_logic ;
  signal R2_PIPE_151_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_5 : std_logic ;
  signal N_5483 : std_logic ;
  signal N_1563 : std_logic ;
  signal R2_PIPE_150_RET : std_logic ;
  signal N_1906 : std_logic ;
  signal R2_PIPE_150_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_6 : std_logic ;
  signal N_5484 : std_logic ;
  signal N_1561 : std_logic ;
  signal R2_PIPE_149_RET : std_logic ;
  signal N_1905 : std_logic ;
  signal R2_PIPE_149_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_7 : std_logic ;
  signal N_5485 : std_logic ;
  signal N_1559 : std_logic ;
  signal R2_PIPE_148_RET : std_logic ;
  signal N_1904 : std_logic ;
  signal R2_PIPE_148_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_8 : std_logic ;
  signal N_5486 : std_logic ;
  signal N_1557 : std_logic ;
  signal R2_PIPE_147_RET : std_logic ;
  signal N_1903 : std_logic ;
  signal R2_PIPE_147_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_9 : std_logic ;
  signal N_5487 : std_logic ;
  signal N_1555 : std_logic ;
  signal R2_PIPE_146_RET : std_logic ;
  signal N_1902 : std_logic ;
  signal R2_PIPE_146_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_10 : std_logic ;
  signal N_5488 : std_logic ;
  signal N_1553 : std_logic ;
  signal R2_PIPE_145_RET : std_logic ;
  signal N_1901 : std_logic ;
  signal R2_PIPE_145_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_11 : std_logic ;
  signal N_5489 : std_logic ;
  signal N_1551 : std_logic ;
  signal R2_PIPE_144_RET : std_logic ;
  signal N_1900 : std_logic ;
  signal R2_PIPE_144_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_12 : std_logic ;
  signal N_5490 : std_logic ;
  signal N_1549 : std_logic ;
  signal R2_PIPE_143_RET : std_logic ;
  signal N_1899 : std_logic ;
  signal R2_PIPE_143_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_13 : std_logic ;
  signal N_5491 : std_logic ;
  signal N_1547 : std_logic ;
  signal R2_PIPE_142_RET : std_logic ;
  signal N_1898 : std_logic ;
  signal R2_PIPE_142_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_14 : std_logic ;
  signal N_5492 : std_logic ;
  signal N_1545 : std_logic ;
  signal R2_PIPE_141_RET : std_logic ;
  signal N_1897 : std_logic ;
  signal R2_PIPE_141_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_15 : std_logic ;
  signal N_5493 : std_logic ;
  signal N_1543 : std_logic ;
  signal R2_PIPE_140_RET : std_logic ;
  signal N_1896 : std_logic ;
  signal R2_PIPE_140_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_16 : std_logic ;
  signal N_5494 : std_logic ;
  signal N_1541 : std_logic ;
  signal R2_PIPE_139_RET : std_logic ;
  signal N_1895 : std_logic ;
  signal R2_PIPE_139_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_17 : std_logic ;
  signal N_5495 : std_logic ;
  signal N_1539 : std_logic ;
  signal R2_PIPE_138_RET : std_logic ;
  signal N_1894 : std_logic ;
  signal R2_PIPE_138_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_18 : std_logic ;
  signal N_5496 : std_logic ;
  signal N_5585 : std_logic ;
  signal N_5586 : std_logic ;
  signal N_5587 : std_logic ;
  signal N_5588 : std_logic ;
  signal N_5589 : std_logic ;
  signal N_5590 : std_logic ;
  signal N_5591 : std_logic ;
  signal N_5592 : std_logic ;
  signal N_5593 : std_logic ;
  signal N_5594 : std_logic ;
  signal N_5595 : std_logic ;
  signal N_5596 : std_logic ;
  signal N_5597 : std_logic ;
  signal N_5598 : std_logic ;
  signal N_5599 : std_logic ;
  signal N_5600 : std_logic ;
  signal N_5601 : std_logic ;
  signal N_5602 : std_logic ;
  signal N_5603 : std_logic ;
  signal N_5604 : std_logic ;
  signal N_5605 : std_logic ;
  signal N_5606 : std_logic ;
  signal N_5607 : std_logic ;
  signal N_5608 : std_logic ;
  signal N_5609 : std_logic ;
  signal N_5610 : std_logic ;
  signal N_5611 : std_logic ;
  signal N_5612 : std_logic ;
  signal N_5613 : std_logic ;
  signal N_5614 : std_logic ;
  signal N_5615 : std_logic ;
  signal N_5616 : std_logic ;
  signal N_5617 : std_logic ;
  signal N_5618 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35 : std_logic ;
  signal R1IN_4_ADD_2_0_CRY_35_RETO_32 : std_logic ;
  signal N_5619 : std_logic ;
  signal UC_187_0 : std_logic ;
  signal UC_188_0 : std_logic ;
  signal UC_189_0 : std_logic ;
  signal UC_190_0 : std_logic ;
  signal UC_191_0 : std_logic ;
  signal UC_192_0 : std_logic ;
  signal UC_193_0 : std_logic ;
  signal UC_194_0 : std_logic ;
  signal UC_195_0 : std_logic ;
  signal UC_196_0 : std_logic ;
  signal UC_197_0 : std_logic ;
  signal UC_198_0 : std_logic ;
  signal UC_199_0 : std_logic ;
  signal UC_200_0 : std_logic ;
  signal UC_173_0 : std_logic ;
  signal UC_174_0 : std_logic ;
  signal UC_175_0 : std_logic ;
  signal UC_176_0 : std_logic ;
  signal UC_177_0 : std_logic ;
  signal UC_178_0 : std_logic ;
  signal UC_179_0 : std_logic ;
  signal UC_180_0 : std_logic ;
  signal UC_181_0 : std_logic ;
  signal UC_182_0 : std_logic ;
  signal UC_183_0 : std_logic ;
  signal UC_184_0 : std_logic ;
  signal UC_185_0 : std_logic ;
  signal UC_186_0 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_1 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_0 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_2 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_1 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_3 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_2 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_4 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_3 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_5 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_4 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_6 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_5 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_7 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_6 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_8 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_7 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_9 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_8 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_10 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_9 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_11 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_10 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_12 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_11 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_13 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_12 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_14 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_13 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_15 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_14 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_16 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_15 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_17 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_16 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_18 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_17 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_19 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_18 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_20 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_19 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_21 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_20 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_22 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_21 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_23 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_22 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_24 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_23 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_25 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_24 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_26 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_25 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_27 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_26 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_28 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_27 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_29 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_28 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_30 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_29 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_31 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_30 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_32 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_31 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_33 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_32 : std_logic ;
  signal R1IN_4_ADD_2_1_0_CRY_33 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_34 : std_logic ;
  signal N_1 : std_logic ;
  signal N_2 : std_logic ;
  signal N_3 : std_logic ;
  signal N_4 : std_logic ;
  signal N_5 : std_logic ;
  signal N_6 : std_logic ;
  signal N_7 : std_logic ;
  signal N_8 : std_logic ;
  signal N_9 : std_logic ;
  signal N_10 : std_logic ;
  signal N_11 : std_logic ;
  signal N_12 : std_logic ;
  signal N_13 : std_logic ;
  signal N_14 : std_logic ;
  signal N_15 : std_logic ;
  signal N_16 : std_logic ;
  signal N_17 : std_logic ;
  signal N_18 : std_logic ;
  signal N_19 : std_logic ;
  signal N_20 : std_logic ;
  signal N_21 : std_logic ;
  signal N_22 : std_logic ;
  signal N_23 : std_logic ;
  signal N_24 : std_logic ;
  signal N_25 : std_logic ;
  signal N_26 : std_logic ;
  signal N_27 : std_logic ;
  signal N_28 : std_logic ;
  signal N_29 : std_logic ;
  signal N_30 : std_logic ;
  signal N_31 : std_logic ;
  signal N_32 : std_logic ;
  signal N_33 : std_logic ;
  signal N_34 : std_logic ;
  signal N_35 : std_logic ;
  signal R2_PIPE_165_RET : std_logic ;
  signal R2_PIPE_165_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_19 : std_logic ;
  signal N_1_0 : std_logic ;
  signal R2_PIPE_164_RET : std_logic ;
  signal R2_PIPE_164_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_20 : std_logic ;
  signal N_1_1 : std_logic ;
  signal R2_PIPE_163_RET : std_logic ;
  signal R2_PIPE_163_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_21 : std_logic ;
  signal N_1_2 : std_logic ;
  signal R2_PIPE_162_RET : std_logic ;
  signal R2_PIPE_162_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_22 : std_logic ;
  signal N_1_3 : std_logic ;
  signal R2_PIPE_161_RET : std_logic ;
  signal R2_PIPE_161_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_23 : std_logic ;
  signal N_1_4 : std_logic ;
  signal R2_PIPE_160_RET : std_logic ;
  signal R2_PIPE_160_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_24 : std_logic ;
  signal N_1_5 : std_logic ;
  signal R2_PIPE_159_RET : std_logic ;
  signal R2_PIPE_159_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_25 : std_logic ;
  signal N_1_6 : std_logic ;
  signal R2_PIPE_158_RET : std_logic ;
  signal R2_PIPE_158_RET_1 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_26 : std_logic ;
  signal N_1_7 : std_logic ;
  signal R1IN_ADD_1_0_CRY_31_RETO_27 : std_logic ;
  signal R1IN_ADD_1_1_0_CRY_28_RETO : std_logic ;
  signal R1IN_ADD_1_1_CRY_28_RETO : std_logic ;
  signal N_1_8 : std_logic ;
  signal N_6019 : std_logic ;
  signal N_6020 : std_logic ;
  signal N_6021 : std_logic ;
  signal N_6022 : std_logic ;
  signal N_6023 : std_logic ;
  signal N_6024 : std_logic ;
  signal N_6025 : std_logic ;
  signal N_6026 : std_logic ;
  signal N_6027 : std_logic ;
  signal N_6028 : std_logic ;
  signal N_6029 : std_logic ;
  signal N_6030 : std_logic ;
  signal N_6031 : std_logic ;
  signal N_6032 : std_logic ;
  signal N_6033 : std_logic ;
  signal N_6034 : std_logic ;
  signal N_6035 : std_logic ;
  signal N_6036 : std_logic ;
  signal N_6037 : std_logic ;
  signal N_6038 : std_logic ;
  signal N_6039 : std_logic ;
  signal N_6040 : std_logic ;
  signal N_6041 : std_logic ;
  signal N_6042 : std_logic ;
  signal N_6043 : std_logic ;
  signal N_6044 : std_logic ;
  signal N_6045 : std_logic ;
  signal N_6046 : std_logic ;
  signal N_6047 : std_logic ;
  signal N_6048 : std_logic ;
  signal N_6049 : std_logic ;
  signal N_6050 : std_logic ;
  signal N_6051 : std_logic ;
  signal N_6052 : std_logic ;
  signal N_6053 : std_logic ;
  signal N_6054 : std_logic ;
  signal N_6055 : std_logic ;
  signal N_6056 : std_logic ;
  signal N_6057 : std_logic ;
  signal N_6058 : std_logic ;
  signal N_6059 : std_logic ;
  signal N_6060 : std_logic ;
  signal N_6061 : std_logic ;
  signal N_1822_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_48 : std_logic ;
  signal N_1821_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_49 : std_logic ;
  signal N_1820_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_93 : std_logic ;
  signal N_1819_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_94 : std_logic ;
  signal N_1818_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_95 : std_logic ;
  signal N_1817_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_96 : std_logic ;
  signal N_1816_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_97 : std_logic ;
  signal N_1815_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_98 : std_logic ;
  signal N_1814_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_99 : std_logic ;
  signal N_1813_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_100 : std_logic ;
  signal N_1812_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_101 : std_logic ;
  signal N_1811_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_102 : std_logic ;
  signal N_1810_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_103 : std_logic ;
  signal N_1809_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_104 : std_logic ;
  signal N_1808_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_105 : std_logic ;
  signal N_1807_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_106 : std_logic ;
  signal N_1806_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_107 : std_logic ;
  signal N_1805_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_108 : std_logic ;
  signal N_1804_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_109 : std_logic ;
  signal N_1803_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_110 : std_logic ;
  signal N_1802_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_111 : std_logic ;
  signal N_1801_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_112 : std_logic ;
  signal N_1800_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_113 : std_logic ;
  signal N_1799_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_114 : std_logic ;
  signal N_1798_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_115 : std_logic ;
  signal N_1797_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_116 : std_logic ;
  signal N_1796_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_117 : std_logic ;
  signal N_1795_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_118 : std_logic ;
  signal N_1794_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_119 : std_logic ;
  signal N_1793_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_120 : std_logic ;
  signal N_1792_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_121 : std_logic ;
  signal N_1791_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_122 : std_logic ;
  signal N_1790_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_123 : std_logic ;
  signal N_1789_RET_0I : std_logic ;
  signal R2_PIPE_104_RET_124 : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_0_RET_0I : std_logic ;
  signal R1IN_4_ADD_2_1_0_AXB_0_RETO : std_logic ;
  signal N_6062 : std_logic ;
  signal N_6402 : std_logic ;
  signal N_6403 : std_logic ;
  signal N_6404 : std_logic ;
  signal N_6405 : std_logic ;
  signal N_6406 : std_logic ;
  signal N_6407 : std_logic ;
  signal N_6408 : std_logic ;
  signal N_6409 : std_logic ;
  signal N_6410 : std_logic ;
  signal N_6411 : std_logic ;
  signal N_6412 : std_logic ;
  signal N_6413 : std_logic ;
  signal N_6414 : std_logic ;
  signal N_6415 : std_logic ;
  signal N_6416 : std_logic ;
  signal N_6417 : std_logic ;
  signal N_6418 : std_logic ;
  signal N_6419 : std_logic ;
  signal N_6420 : std_logic ;
  signal N_6421 : std_logic ;
  signal N_6422 : std_logic ;
  signal N_6423 : std_logic ;
  signal N_6424 : std_logic ;
  signal N_6425 : std_logic ;
  signal N_6426 : std_logic ;
  signal N_6427 : std_logic ;
  signal N_6428 : std_logic ;
  signal N_6429 : std_logic ;
  signal N_6430 : std_logic ;
  signal N_6431 : std_logic ;
  signal N_6432 : std_logic ;
  signal N_6433 : std_logic ;
  signal N_6434 : std_logic ;
  signal N_6435 : std_logic ;
  signal N_6436 : std_logic ;
  signal N_6437 : std_logic ;
  signal N_6438 : std_logic ;
  signal N_6439 : std_logic ;
  signal N_6440 : std_logic ;
  signal N_6441 : std_logic ;
  signal N_6442 : std_logic ;
  signal N_6443 : std_logic ;
  signal N_6444 : std_logic ;
  signal N_6445 : std_logic ;
  signal N_6446 : std_logic ;
  signal N_6447 : std_logic ;
  signal N_6448 : std_logic ;
  signal N_6449 : std_logic ;
  signal N_6450 : std_logic ;
  signal N_6451 : std_logic ;
  signal N_6452 : std_logic ;
  signal N_6453 : std_logic ;
  signal N_6454 : std_logic ;
  signal N_6455 : std_logic ;
  signal N_6456 : std_logic ;
  signal N_6457 : std_logic ;
  signal N_6458 : std_logic ;
  signal N_6459 : std_logic ;
  signal N_6460 : std_logic ;
  signal N_6461 : std_logic ;
  signal N_6462 : std_logic ;
  signal N_6463 : std_logic ;
  signal N_6464 : std_logic ;
  signal N_6465 : std_logic ;
  signal N_6466 : std_logic ;
  signal N_6467 : std_logic ;
  signal N_6468 : std_logic ;
  signal N_6469 : std_logic ;
  signal N_6470 : std_logic ;
  signal N_6471 : std_logic ;
  signal N_6472 : std_logic ;
  signal N_6473 : std_logic ;
  signal N_6474 : std_logic ;
  signal N_6475 : std_logic ;
  signal N_6476 : std_logic ;
  signal N_6477 : std_logic ;
  signal N_6478 : std_logic ;
  signal N_6479 : std_logic ;
  signal N_6480 : std_logic ;
  signal N_6654 : std_logic ;
  signal N_6655 : std_logic ;
  signal N_6656 : std_logic ;
  signal N_6657 : std_logic ;
  signal N_6658 : std_logic ;
  signal N_6659 : std_logic ;
  signal N_6660 : std_logic ;
  signal N_6661 : std_logic ;
  signal N_6662 : std_logic ;
  signal N_6663 : std_logic ;
  signal N_6664 : std_logic ;
  signal N_6665 : std_logic ;
  signal N_6666 : std_logic ;
  signal N_6667 : std_logic ;
  signal N_6668 : std_logic ;
  signal N_6669 : std_logic ;
  signal N_6670 : std_logic ;
  signal N_6671 : std_logic ;
  signal N_6672 : std_logic ;
  signal N_6673 : std_logic ;
  signal N_6674 : std_logic ;
  signal N_6675 : std_logic ;
  signal N_6676 : std_logic ;
  signal N_6677 : std_logic ;
  signal N_6678 : std_logic ;
  signal N_6679 : std_logic ;
  signal N_6680 : std_logic ;
  signal N_6681 : std_logic ;
  signal N_6682 : std_logic ;
  signal N_6683 : std_logic ;
  signal N_6684 : std_logic ;
  signal N_6685 : std_logic ;
  signal N_6686 : std_logic ;
  signal N_6687 : std_logic ;
  signal N_6688 : std_logic ;
  signal N_6689 : std_logic ;
  signal N_6690 : std_logic ;
  signal N_6691 : std_logic ;
  signal N_6692 : std_logic ;
  signal N_6693 : std_logic ;
  signal N_6694 : std_logic ;
  signal N_6695 : std_logic ;
  signal N_6696 : std_logic ;
  signal N_6697 : std_logic ;
  signal N_6698 : std_logic ;
  signal N_6699 : std_logic ;
  signal N_6700 : std_logic ;
  signal N_6701 : std_logic ;
  signal N_6702 : std_logic ;
  signal N_6703 : std_logic ;
  signal N_6704 : std_logic ;
  signal N_6705 : std_logic ;
  signal N_6706 : std_logic ;
  signal N_6707 : std_logic ;
  signal N_6708 : std_logic ;
  signal N_6709 : std_logic ;
  signal N_6710 : std_logic ;
  signal N_6711 : std_logic ;
  signal N_6712 : std_logic ;
  signal N_6713 : std_logic ;
  signal N_6714 : std_logic ;
  signal N_6715 : std_logic ;
  signal N_6716 : std_logic ;
  signal N_6717 : std_logic ;
  signal N_6718 : std_logic ;
  signal N_6719 : std_logic ;
  signal N_6720 : std_logic ;
  signal N_6721 : std_logic ;
  signal N_6722 : std_logic ;
  signal N_6723 : std_logic ;
  signal N_6724 : std_logic ;
  signal N_6725 : std_logic ;
  signal N_6726 : std_logic ;
  signal N_6727 : std_logic ;
  signal N_6728 : std_logic ;
  signal N_6729 : std_logic ;
  signal N_6730 : std_logic ;
  signal N_6731 : std_logic ;
  signal N_6732 : std_logic ;
  signal N_6906 : std_logic ;
  signal N_6907 : std_logic ;
  signal N_6908 : std_logic ;
  signal N_6909 : std_logic ;
  signal N_6910 : std_logic ;
  signal N_6911 : std_logic ;
  signal N_6912 : std_logic ;
  signal N_6913 : std_logic ;
  signal N_6914 : std_logic ;
  signal N_6915 : std_logic ;
  signal N_6916 : std_logic ;
  signal N_6917 : std_logic ;
  signal N_6918 : std_logic ;
  signal N_6919 : std_logic ;
  signal N_6920 : std_logic ;
  signal N_6921 : std_logic ;
  signal N_6922 : std_logic ;
  signal N_6923 : std_logic ;
  signal N_6924 : std_logic ;
  signal N_6925 : std_logic ;
  signal N_6926 : std_logic ;
  signal N_6927 : std_logic ;
  signal N_6928 : std_logic ;
  signal N_6929 : std_logic ;
  signal N_6930 : std_logic ;
  signal N_6931 : std_logic ;
  signal N_6932 : std_logic ;
  signal N_6933 : std_logic ;
  signal N_6934 : std_logic ;
  signal N_6935 : std_logic ;
  signal N_6936 : std_logic ;
  signal N_6937 : std_logic ;
  signal N_6938 : std_logic ;
  signal N_6939 : std_logic ;
  signal N_6940 : std_logic ;
  signal N_6941 : std_logic ;
  signal N_6942 : std_logic ;
  signal N_6943 : std_logic ;
  signal N_6944 : std_logic ;
  signal N_6945 : std_logic ;
  signal N_6946 : std_logic ;
  signal N_6947 : std_logic ;
  signal N_6948 : std_logic ;
  signal N_6949 : std_logic ;
  signal N_6950 : std_logic ;
  signal N_6951 : std_logic ;
  signal N_6952 : std_logic ;
  signal N_6953 : std_logic ;
  signal N_6954 : std_logic ;
  signal N_6955 : std_logic ;
  signal N_6956 : std_logic ;
  signal N_6957 : std_logic ;
  signal N_6958 : std_logic ;
  signal N_6959 : std_logic ;
  signal N_6960 : std_logic ;
  signal N_6961 : std_logic ;
  signal N_6962 : std_logic ;
  signal N_6963 : std_logic ;
  signal N_6964 : std_logic ;
  signal N_6965 : std_logic ;
  signal N_6966 : std_logic ;
  signal N_6967 : std_logic ;
  signal N_6968 : std_logic ;
  signal N_6969 : std_logic ;
  signal N_6970 : std_logic ;
  signal N_6971 : std_logic ;
  signal N_6972 : std_logic ;
  signal N_6973 : std_logic ;
  signal N_6974 : std_logic ;
  signal N_6975 : std_logic ;
  signal N_6976 : std_logic ;
  signal N_6977 : std_logic ;
  signal N_6978 : std_logic ;
  signal N_6979 : std_logic ;
  signal N_6980 : std_logic ;
  signal N_6981 : std_logic ;
  signal N_6982 : std_logic ;
  signal N_6983 : std_logic ;
  signal N_6984 : std_logic ;
  signal N_7158 : std_logic ;
  signal N_7159 : std_logic ;
  signal N_7160 : std_logic ;
  signal N_7161 : std_logic ;
  signal N_7162 : std_logic ;
  signal N_7163 : std_logic ;
  signal N_7164 : std_logic ;
  signal N_7165 : std_logic ;
  signal N_7166 : std_logic ;
  signal N_7167 : std_logic ;
  signal N_7168 : std_logic ;
  signal N_7169 : std_logic ;
  signal N_7170 : std_logic ;
  signal N_7171 : std_logic ;
  signal N_7172 : std_logic ;
  signal N_7173 : std_logic ;
  signal N_7174 : std_logic ;
  signal N_7175 : std_logic ;
  signal N_7176 : std_logic ;
  signal N_7177 : std_logic ;
  signal N_7178 : std_logic ;
  signal N_7179 : std_logic ;
  signal N_7180 : std_logic ;
  signal N_7181 : std_logic ;
  signal N_7182 : std_logic ;
  signal N_7183 : std_logic ;
  signal N_7184 : std_logic ;
  signal N_7185 : std_logic ;
  signal N_7186 : std_logic ;
  signal N_7187 : std_logic ;
  signal N_7188 : std_logic ;
  signal N_7189 : std_logic ;
  signal N_7190 : std_logic ;
  signal N_7191 : std_logic ;
  signal N_7192 : std_logic ;
  signal N_7193 : std_logic ;
  signal N_7194 : std_logic ;
  signal N_7195 : std_logic ;
  signal N_7196 : std_logic ;
  signal N_7197 : std_logic ;
  signal N_7198 : std_logic ;
  signal N_7199 : std_logic ;
  signal N_7200 : std_logic ;
  signal N_7201 : std_logic ;
  signal N_7202 : std_logic ;
  signal N_7203 : std_logic ;
  signal N_7204 : std_logic ;
  signal N_7205 : std_logic ;
  signal N_7206 : std_logic ;
  signal N_7207 : std_logic ;
  signal N_7208 : std_logic ;
  signal N_7209 : std_logic ;
  signal N_7210 : std_logic ;
  signal N_7211 : std_logic ;
  signal N_7212 : std_logic ;
  signal N_7213 : std_logic ;
  signal N_7214 : std_logic ;
  signal N_7215 : std_logic ;
  signal N_7216 : std_logic ;
  signal N_7217 : std_logic ;
  signal N_7218 : std_logic ;
  signal N_7219 : std_logic ;
  signal N_7220 : std_logic ;
  signal N_7221 : std_logic ;
  signal N_7222 : std_logic ;
  signal N_7223 : std_logic ;
  signal N_7224 : std_logic ;
  signal N_7225 : std_logic ;
  signal N_7226 : std_logic ;
  signal N_7227 : std_logic ;
  signal N_7228 : std_logic ;
  signal N_7229 : std_logic ;
  signal N_7230 : std_logic ;
  signal N_7231 : std_logic ;
  signal N_7232 : std_logic ;
  signal N_7233 : std_logic ;
  signal N_7234 : std_logic ;
  signal N_7235 : std_logic ;
  signal N_7236 : std_logic ;
  signal N_7410 : std_logic ;
  signal N_7411 : std_logic ;
  signal N_7412 : std_logic ;
  signal N_7413 : std_logic ;
  signal N_7414 : std_logic ;
  signal N_7415 : std_logic ;
  signal N_7416 : std_logic ;
  signal N_7417 : std_logic ;
  signal N_7418 : std_logic ;
  signal N_7419 : std_logic ;
  signal N_7420 : std_logic ;
  signal N_7421 : std_logic ;
  signal N_7422 : std_logic ;
  signal N_7423 : std_logic ;
  signal N_7424 : std_logic ;
  signal N_7425 : std_logic ;
  signal N_7426 : std_logic ;
  signal N_7427 : std_logic ;
  signal N_7428 : std_logic ;
  signal N_7429 : std_logic ;
  signal N_7430 : std_logic ;
  signal N_7431 : std_logic ;
  signal N_7432 : std_logic ;
  signal N_7433 : std_logic ;
  signal N_7434 : std_logic ;
  signal N_7435 : std_logic ;
  signal N_7436 : std_logic ;
  signal N_7437 : std_logic ;
  signal N_7438 : std_logic ;
  signal N_7439 : std_logic ;
  signal N_7440 : std_logic ;
  signal N_7441 : std_logic ;
  signal N_7442 : std_logic ;
  signal N_7443 : std_logic ;
  signal N_7444 : std_logic ;
  signal N_7445 : std_logic ;
  signal N_7446 : std_logic ;
  signal N_7447 : std_logic ;
  signal N_7448 : std_logic ;
  signal N_7449 : std_logic ;
  signal N_7450 : std_logic ;
  signal N_7451 : std_logic ;
  signal N_7452 : std_logic ;
  signal N_7453 : std_logic ;
  signal N_7454 : std_logic ;
  signal N_7455 : std_logic ;
  signal N_7456 : std_logic ;
  signal N_7457 : std_logic ;
  signal N_7458 : std_logic ;
  signal N_7459 : std_logic ;
  signal N_7460 : std_logic ;
  signal N_7461 : std_logic ;
  signal N_7462 : std_logic ;
  signal N_7463 : std_logic ;
  signal N_7464 : std_logic ;
  signal N_7465 : std_logic ;
  signal N_7466 : std_logic ;
  signal N_7467 : std_logic ;
  signal N_7468 : std_logic ;
  signal N_7469 : std_logic ;
  signal N_7470 : std_logic ;
  signal N_7471 : std_logic ;
  signal N_7472 : std_logic ;
  signal N_7473 : std_logic ;
  signal N_7474 : std_logic ;
  signal N_7475 : std_logic ;
  signal N_7476 : std_logic ;
  signal N_7477 : std_logic ;
  signal N_7478 : std_logic ;
  signal N_7479 : std_logic ;
  signal N_7480 : std_logic ;
  signal N_7481 : std_logic ;
  signal N_7482 : std_logic ;
  signal N_7483 : std_logic ;
  signal N_7484 : std_logic ;
  signal N_7485 : std_logic ;
  signal N_7486 : std_logic ;
  signal N_7487 : std_logic ;
  signal N_7488 : std_logic ;
  signal N_8038 : std_logic ;
  signal N_8039 : std_logic ;
  signal N_8040 : std_logic ;
  signal N_8041 : std_logic ;
  signal N_8042 : std_logic ;
  signal N_8043 : std_logic ;
  signal N_8044 : std_logic ;
  signal N_8045 : std_logic ;
  signal N_8046 : std_logic ;
  signal N_8047 : std_logic ;
  signal N_8048 : std_logic ;
  signal N_8049 : std_logic ;
  signal N_8050 : std_logic ;
  signal N_8051 : std_logic ;
  signal N_8052 : std_logic ;
  signal N_8053 : std_logic ;
  signal N_8054 : std_logic ;
  signal N_8055 : std_logic ;
  signal N_8056 : std_logic ;
  signal N_8057 : std_logic ;
  signal N_8058 : std_logic ;
  signal N_8059 : std_logic ;
  signal N_8060 : std_logic ;
  signal N_8061 : std_logic ;
  signal N_8062 : std_logic ;
  signal N_8063 : std_logic ;
  signal N_8064 : std_logic ;
  signal N_8065 : std_logic ;
  signal N_8066 : std_logic ;
  signal N_8067 : std_logic ;
  signal N_8068 : std_logic ;
  signal N_8069 : std_logic ;
  signal N_8070 : std_logic ;
  signal N_8071 : std_logic ;
  signal N_8072 : std_logic ;
  signal N_8073 : std_logic ;
  signal N_8074 : std_logic ;
  signal N_8075 : std_logic ;
  signal N_8076 : std_logic ;
  signal N_8077 : std_logic ;
  signal N_8078 : std_logic ;
  signal N_8079 : std_logic ;
  signal N_8080 : std_logic ;
  signal N_8081 : std_logic ;
  signal N_8082 : std_logic ;
  signal N_8083 : std_logic ;
  signal N_8084 : std_logic ;
  signal N_8085 : std_logic ;
  signal N_8086 : std_logic ;
  signal N_8087 : std_logic ;
  signal N_8088 : std_logic ;
  signal N_8089 : std_logic ;
  signal N_8090 : std_logic ;
  signal N_8091 : std_logic ;
  signal N_8092 : std_logic ;
  signal N_8093 : std_logic ;
  signal N_8094 : std_logic ;
  signal N_8095 : std_logic ;
  signal N_8096 : std_logic ;
  signal N_8097 : std_logic ;
  signal N_8098 : std_logic ;
  signal N_8099 : std_logic ;
  signal N_8100 : std_logic ;
  signal N_8101 : std_logic ;
  signal N_8102 : std_logic ;
  signal N_8103 : std_logic ;
  signal N_8104 : std_logic ;
  signal N_8105 : std_logic ;
  signal N_8106 : std_logic ;
  signal N_8107 : std_logic ;
  signal N_8108 : std_logic ;
  signal N_8109 : std_logic ;
  signal N_8110 : std_logic ;
  signal N_8111 : std_logic ;
  signal N_8112 : std_logic ;
  signal N_8113 : std_logic ;
  signal N_8114 : std_logic ;
  signal N_8115 : std_logic ;
  signal N_8116 : std_logic ;
  signal N_8290 : std_logic ;
  signal N_8291 : std_logic ;
  signal N_8292 : std_logic ;
  signal N_8293 : std_logic ;
  signal N_8294 : std_logic ;
  signal N_8295 : std_logic ;
  signal N_8296 : std_logic ;
  signal N_8297 : std_logic ;
  signal N_8298 : std_logic ;
  signal N_8299 : std_logic ;
  signal N_8300 : std_logic ;
  signal N_8301 : std_logic ;
  signal N_8302 : std_logic ;
  signal N_8303 : std_logic ;
  signal N_8304 : std_logic ;
  signal N_8305 : std_logic ;
  signal N_8306 : std_logic ;
  signal N_8307 : std_logic ;
  signal N_8308 : std_logic ;
  signal N_8309 : std_logic ;
  signal N_8310 : std_logic ;
  signal N_8311 : std_logic ;
  signal N_8312 : std_logic ;
  signal N_8313 : std_logic ;
  signal N_8314 : std_logic ;
  signal N_8315 : std_logic ;
  signal N_8316 : std_logic ;
  signal N_8317 : std_logic ;
  signal N_8318 : std_logic ;
  signal N_8319 : std_logic ;
  signal N_8320 : std_logic ;
  signal N_8321 : std_logic ;
  signal N_8322 : std_logic ;
  signal N_8323 : std_logic ;
  signal N_8324 : std_logic ;
  signal N_8325 : std_logic ;
  signal N_8326 : std_logic ;
  signal N_8327 : std_logic ;
  signal N_8328 : std_logic ;
  signal N_8329 : std_logic ;
  signal N_8330 : std_logic ;
  signal N_8331 : std_logic ;
  signal N_8332 : std_logic ;
  signal N_8333 : std_logic ;
  signal N_8334 : std_logic ;
  signal N_8335 : std_logic ;
  signal N_8336 : std_logic ;
  signal N_8337 : std_logic ;
  signal N_8338 : std_logic ;
  signal N_8339 : std_logic ;
  signal N_8340 : std_logic ;
  signal N_8341 : std_logic ;
  signal N_8342 : std_logic ;
  signal N_8343 : std_logic ;
  signal N_8344 : std_logic ;
  signal N_8345 : std_logic ;
  signal N_8346 : std_logic ;
  signal N_8347 : std_logic ;
  signal N_8348 : std_logic ;
  signal N_8349 : std_logic ;
  signal N_8350 : std_logic ;
  signal N_8351 : std_logic ;
  signal N_8352 : std_logic ;
  signal N_8353 : std_logic ;
  signal N_8354 : std_logic ;
  signal N_8355 : std_logic ;
  signal N_8356 : std_logic ;
  signal N_8357 : std_logic ;
  signal N_8358 : std_logic ;
  signal N_8359 : std_logic ;
  signal N_8360 : std_logic ;
  signal N_8361 : std_logic ;
  signal N_8362 : std_logic ;
  signal N_8363 : std_logic ;
  signal N_8364 : std_logic ;
  signal N_8365 : std_logic ;
  signal N_8366 : std_logic ;
  signal N_8367 : std_logic ;
  signal N_8368 : std_logic ;
  signal N_8542 : std_logic ;
  signal N_8543 : std_logic ;
  signal N_8544 : std_logic ;
  signal N_8545 : std_logic ;
  signal N_8546 : std_logic ;
  signal N_8547 : std_logic ;
  signal N_8548 : std_logic ;
  signal N_8549 : std_logic ;
  signal N_8550 : std_logic ;
  signal N_8551 : std_logic ;
  signal N_8552 : std_logic ;
  signal N_8553 : std_logic ;
  signal N_8554 : std_logic ;
  signal N_8555 : std_logic ;
  signal N_8556 : std_logic ;
  signal N_8557 : std_logic ;
  signal N_8558 : std_logic ;
  signal N_8559 : std_logic ;
  signal N_8560 : std_logic ;
  signal N_8561 : std_logic ;
  signal N_8562 : std_logic ;
  signal N_8563 : std_logic ;
  signal N_8564 : std_logic ;
  signal N_8565 : std_logic ;
  signal N_8566 : std_logic ;
  signal N_8567 : std_logic ;
  signal N_8568 : std_logic ;
  signal N_8569 : std_logic ;
  signal N_8570 : std_logic ;
  signal N_8571 : std_logic ;
  signal N_8572 : std_logic ;
  signal N_8573 : std_logic ;
  signal N_8574 : std_logic ;
  signal N_8575 : std_logic ;
  signal N_8576 : std_logic ;
  signal N_8577 : std_logic ;
  signal N_8578 : std_logic ;
  signal N_8579 : std_logic ;
  signal N_8580 : std_logic ;
  signal N_8581 : std_logic ;
  signal N_8582 : std_logic ;
  signal N_8583 : std_logic ;
  signal N_8584 : std_logic ;
  signal N_8585 : std_logic ;
  signal N_8586 : std_logic ;
  signal N_8587 : std_logic ;
  signal N_8588 : std_logic ;
  signal N_8589 : std_logic ;
  signal N_8590 : std_logic ;
  signal N_8591 : std_logic ;
  signal N_8592 : std_logic ;
  signal N_8593 : std_logic ;
  signal N_8594 : std_logic ;
  signal N_8595 : std_logic ;
  signal N_8596 : std_logic ;
  signal N_8597 : std_logic ;
  signal N_8598 : std_logic ;
  signal N_8599 : std_logic ;
  signal N_8600 : std_logic ;
  signal N_8601 : std_logic ;
  signal N_8602 : std_logic ;
  signal N_8603 : std_logic ;
  signal N_8604 : std_logic ;
  signal N_8605 : std_logic ;
  signal N_8606 : std_logic ;
  signal N_8607 : std_logic ;
  signal N_8608 : std_logic ;
  signal N_8609 : std_logic ;
  signal N_8610 : std_logic ;
  signal N_8611 : std_logic ;
  signal N_8612 : std_logic ;
  signal N_8613 : std_logic ;
  signal N_8614 : std_logic ;
  signal N_8615 : std_logic ;
  signal N_8616 : std_logic ;
  signal N_8617 : std_logic ;
  signal N_8618 : std_logic ;
  signal N_8619 : std_logic ;
  signal N_8620 : std_logic ;
  signal N_9170 : std_logic ;
  signal N_9171 : std_logic ;
  signal N_9172 : std_logic ;
  signal N_9173 : std_logic ;
  signal N_9174 : std_logic ;
  signal N_9175 : std_logic ;
  signal N_9176 : std_logic ;
  signal N_9177 : std_logic ;
  signal N_9178 : std_logic ;
  signal N_9179 : std_logic ;
  signal N_9180 : std_logic ;
  signal N_9181 : std_logic ;
  signal N_9182 : std_logic ;
  signal N_9183 : std_logic ;
  signal N_9184 : std_logic ;
  signal N_9185 : std_logic ;
  signal N_9186 : std_logic ;
  signal N_9187 : std_logic ;
  signal N_9188 : std_logic ;
  signal N_9189 : std_logic ;
  signal N_9190 : std_logic ;
  signal N_9191 : std_logic ;
  signal N_9192 : std_logic ;
  signal N_9193 : std_logic ;
  signal N_9194 : std_logic ;
  signal N_9195 : std_logic ;
  signal N_9196 : std_logic ;
  signal N_9197 : std_logic ;
  signal N_9198 : std_logic ;
  signal N_9199 : std_logic ;
  signal N_9200 : std_logic ;
  signal N_9201 : std_logic ;
  signal N_9202 : std_logic ;
  signal N_9203 : std_logic ;
  signal N_9204 : std_logic ;
  signal N_9205 : std_logic ;
  signal N_9206 : std_logic ;
  signal N_9207 : std_logic ;
  signal N_9208 : std_logic ;
  signal N_9209 : std_logic ;
  signal N_9210 : std_logic ;
  signal N_9211 : std_logic ;
  signal N_9212 : std_logic ;
  signal N_9213 : std_logic ;
  signal N_9214 : std_logic ;
  signal N_9215 : std_logic ;
  signal N_9216 : std_logic ;
  signal N_9217 : std_logic ;
  signal N_9218 : std_logic ;
  signal N_9219 : std_logic ;
  signal N_9220 : std_logic ;
  signal N_9221 : std_logic ;
  signal N_9222 : std_logic ;
  signal N_9223 : std_logic ;
  signal N_9224 : std_logic ;
  signal N_9225 : std_logic ;
  signal N_9226 : std_logic ;
  signal N_9227 : std_logic ;
  signal N_9228 : std_logic ;
  signal N_9229 : std_logic ;
  signal N_9230 : std_logic ;
  signal N_9231 : std_logic ;
  signal N_9232 : std_logic ;
  signal N_9233 : std_logic ;
  signal N_9234 : std_logic ;
  signal N_9235 : std_logic ;
  signal N_9236 : std_logic ;
  signal N_9237 : std_logic ;
  signal N_9238 : std_logic ;
  signal N_9239 : std_logic ;
  signal N_9240 : std_logic ;
  signal N_9241 : std_logic ;
  signal N_9242 : std_logic ;
  signal N_9243 : std_logic ;
  signal N_9244 : std_logic ;
  signal N_9245 : std_logic ;
  signal N_9246 : std_logic ;
  signal N_9247 : std_logic ;
  signal N_9248 : std_logic ;
  signal N_9422 : std_logic ;
  signal N_9423 : std_logic ;
  signal N_9424 : std_logic ;
  signal N_9425 : std_logic ;
  signal N_9426 : std_logic ;
  signal N_9427 : std_logic ;
  signal N_9428 : std_logic ;
  signal N_9429 : std_logic ;
  signal N_9430 : std_logic ;
  signal N_9431 : std_logic ;
  signal N_9432 : std_logic ;
  signal N_9433 : std_logic ;
  signal N_9434 : std_logic ;
  signal N_9435 : std_logic ;
  signal N_9436 : std_logic ;
  signal N_9437 : std_logic ;
  signal N_9438 : std_logic ;
  signal N_9439 : std_logic ;
  signal N_9440 : std_logic ;
  signal N_9441 : std_logic ;
  signal N_9442 : std_logic ;
  signal N_9443 : std_logic ;
  signal N_9444 : std_logic ;
  signal N_9445 : std_logic ;
  signal N_9446 : std_logic ;
  signal N_9447 : std_logic ;
  signal N_9448 : std_logic ;
  signal N_9449 : std_logic ;
  signal N_9450 : std_logic ;
  signal N_9451 : std_logic ;
  signal N_9452 : std_logic ;
  signal N_9453 : std_logic ;
  signal N_9454 : std_logic ;
  signal N_9455 : std_logic ;
  signal N_9456 : std_logic ;
  signal N_9457 : std_logic ;
  signal N_9458 : std_logic ;
  signal N_9459 : std_logic ;
  signal N_9460 : std_logic ;
  signal N_9461 : std_logic ;
  signal N_9462 : std_logic ;
  signal N_9463 : std_logic ;
  signal N_9464 : std_logic ;
  signal N_9465 : std_logic ;
  signal N_9466 : std_logic ;
  signal N_9467 : std_logic ;
  signal N_9468 : std_logic ;
  signal N_9469 : std_logic ;
  signal N_9470 : std_logic ;
  signal N_9471 : std_logic ;
  signal N_9472 : std_logic ;
  signal N_9473 : std_logic ;
  signal N_9474 : std_logic ;
  signal N_9475 : std_logic ;
  signal N_9476 : std_logic ;
  signal N_9477 : std_logic ;
  signal N_9478 : std_logic ;
  signal N_9479 : std_logic ;
  signal N_9480 : std_logic ;
  signal N_9481 : std_logic ;
  signal N_9482 : std_logic ;
  signal N_9483 : std_logic ;
  signal N_9484 : std_logic ;
  signal N_9485 : std_logic ;
  signal N_9486 : std_logic ;
  signal N_9487 : std_logic ;
  signal N_9488 : std_logic ;
  signal N_9489 : std_logic ;
  signal N_9490 : std_logic ;
  signal N_9491 : std_logic ;
  signal N_9492 : std_logic ;
  signal N_9493 : std_logic ;
  signal N_9494 : std_logic ;
  signal N_9495 : std_logic ;
  signal N_9496 : std_logic ;
  signal N_9497 : std_logic ;
  signal N_9498 : std_logic ;
  signal N_9499 : std_logic ;
  signal N_9500 : std_logic ;
  signal N_9674 : std_logic ;
  signal N_9675 : std_logic ;
  signal N_9676 : std_logic ;
  signal N_9677 : std_logic ;
  signal N_9678 : std_logic ;
  signal N_9679 : std_logic ;
  signal N_9680 : std_logic ;
  signal N_9681 : std_logic ;
  signal N_9682 : std_logic ;
  signal N_9683 : std_logic ;
  signal N_9684 : std_logic ;
  signal N_9685 : std_logic ;
  signal N_9686 : std_logic ;
  signal N_9687 : std_logic ;
  signal N_9688 : std_logic ;
  signal N_9689 : std_logic ;
  signal N_9690 : std_logic ;
  signal N_9691 : std_logic ;
  signal N_9692 : std_logic ;
  signal N_9693 : std_logic ;
  signal N_9694 : std_logic ;
  signal N_9695 : std_logic ;
  signal N_9696 : std_logic ;
  signal N_9697 : std_logic ;
  signal N_9698 : std_logic ;
  signal N_9699 : std_logic ;
  signal N_9700 : std_logic ;
  signal N_9701 : std_logic ;
  signal N_9702 : std_logic ;
  signal N_9703 : std_logic ;
  signal N_9704 : std_logic ;
  signal N_9705 : std_logic ;
  signal N_9706 : std_logic ;
  signal N_9707 : std_logic ;
  signal N_9708 : std_logic ;
  signal N_9709 : std_logic ;
  signal N_9710 : std_logic ;
  signal N_9711 : std_logic ;
  signal N_9712 : std_logic ;
  signal N_9713 : std_logic ;
  signal N_9714 : std_logic ;
  signal N_9715 : std_logic ;
  signal N_9716 : std_logic ;
  signal N_9717 : std_logic ;
  signal N_9718 : std_logic ;
  signal N_9719 : std_logic ;
  signal N_9720 : std_logic ;
  signal N_9721 : std_logic ;
  signal N_9722 : std_logic ;
  signal N_9723 : std_logic ;
  signal N_9724 : std_logic ;
  signal N_9725 : std_logic ;
  signal N_9726 : std_logic ;
  signal N_9727 : std_logic ;
  signal N_9728 : std_logic ;
  signal N_9729 : std_logic ;
  signal N_9730 : std_logic ;
  signal N_9731 : std_logic ;
  signal N_9732 : std_logic ;
  signal N_9733 : std_logic ;
  signal N_9734 : std_logic ;
  signal N_9735 : std_logic ;
  signal N_9736 : std_logic ;
  signal N_9737 : std_logic ;
  signal N_9738 : std_logic ;
  signal N_9739 : std_logic ;
  signal N_9740 : std_logic ;
  signal N_9741 : std_logic ;
  signal N_9742 : std_logic ;
  signal N_9743 : std_logic ;
  signal N_9744 : std_logic ;
  signal N_9745 : std_logic ;
  signal N_9746 : std_logic ;
  signal N_9747 : std_logic ;
  signal N_9748 : std_logic ;
  signal N_9749 : std_logic ;
  signal N_9750 : std_logic ;
  signal N_9751 : std_logic ;
  signal N_9752 : std_logic ;
  signal N_10302 : std_logic ;
  signal N_10303 : std_logic ;
  signal N_10304 : std_logic ;
  signal N_10305 : std_logic ;
  signal N_10306 : std_logic ;
  signal N_10307 : std_logic ;
  signal N_10308 : std_logic ;
  signal N_10309 : std_logic ;
  signal N_10310 : std_logic ;
  signal N_10311 : std_logic ;
  signal N_10312 : std_logic ;
  signal N_10313 : std_logic ;
  signal N_10314 : std_logic ;
  signal N_10315 : std_logic ;
  signal N_10316 : std_logic ;
  signal N_10317 : std_logic ;
  signal N_10318 : std_logic ;
  signal N_10319 : std_logic ;
  signal N_10320 : std_logic ;
  signal N_10321 : std_logic ;
  signal N_10322 : std_logic ;
  signal N_10323 : std_logic ;
  signal N_10324 : std_logic ;
  signal N_10325 : std_logic ;
  signal N_10326 : std_logic ;
  signal N_10327 : std_logic ;
  signal N_10328 : std_logic ;
  signal N_10329 : std_logic ;
  signal N_10330 : std_logic ;
  signal N_10331 : std_logic ;
  signal N_10332 : std_logic ;
  signal N_10333 : std_logic ;
  signal N_10334 : std_logic ;
  signal N_10335 : std_logic ;
  signal N_10336 : std_logic ;
  signal N_10337 : std_logic ;
  signal N_10338 : std_logic ;
  signal N_10339 : std_logic ;
  signal N_10340 : std_logic ;
  signal N_10341 : std_logic ;
  signal N_10342 : std_logic ;
  signal N_10343 : std_logic ;
  signal N_10344 : std_logic ;
  signal N_10345 : std_logic ;
  signal N_10346 : std_logic ;
  signal N_10347 : std_logic ;
  signal N_10348 : std_logic ;
  signal N_10349 : std_logic ;
  signal N_10350 : std_logic ;
  signal N_10351 : std_logic ;
  signal N_10352 : std_logic ;
  signal N_10353 : std_logic ;
  signal N_10354 : std_logic ;
  signal N_10355 : std_logic ;
  signal N_10356 : std_logic ;
  signal N_10357 : std_logic ;
  signal N_10358 : std_logic ;
  signal N_10359 : std_logic ;
  signal N_10360 : std_logic ;
  signal N_10361 : std_logic ;
  signal N_10362 : std_logic ;
  signal N_10363 : std_logic ;
  signal N_10364 : std_logic ;
  signal N_10365 : std_logic ;
  signal N_10366 : std_logic ;
  signal N_10367 : std_logic ;
  signal N_10368 : std_logic ;
  signal N_10369 : std_logic ;
  signal N_10370 : std_logic ;
  signal N_10371 : std_logic ;
  signal N_10372 : std_logic ;
  signal N_10373 : std_logic ;
  signal N_10374 : std_logic ;
  signal N_10375 : std_logic ;
  signal N_10376 : std_logic ;
  signal N_10377 : std_logic ;
  signal N_10378 : std_logic ;
  signal N_10379 : std_logic ;
  signal N_10380 : std_logic ;
  signal N_10554 : std_logic ;
  signal N_10555 : std_logic ;
  signal N_10556 : std_logic ;
  signal N_10557 : std_logic ;
  signal N_10558 : std_logic ;
  signal N_10559 : std_logic ;
  signal N_10560 : std_logic ;
  signal N_10561 : std_logic ;
  signal N_10562 : std_logic ;
  signal N_10563 : std_logic ;
  signal N_10564 : std_logic ;
  signal N_10565 : std_logic ;
  signal N_10566 : std_logic ;
  signal N_10567 : std_logic ;
  signal N_10568 : std_logic ;
  signal N_10569 : std_logic ;
  signal N_10570 : std_logic ;
  signal N_10571 : std_logic ;
  signal N_10572 : std_logic ;
  signal N_10573 : std_logic ;
  signal N_10574 : std_logic ;
  signal N_10575 : std_logic ;
  signal N_10576 : std_logic ;
  signal N_10577 : std_logic ;
  signal N_10578 : std_logic ;
  signal N_10579 : std_logic ;
  signal N_10580 : std_logic ;
  signal N_10581 : std_logic ;
  signal N_10582 : std_logic ;
  signal N_10583 : std_logic ;
  signal N_10584 : std_logic ;
  signal N_10585 : std_logic ;
  signal N_10586 : std_logic ;
  signal N_10587 : std_logic ;
  signal N_10588 : std_logic ;
  signal N_10589 : std_logic ;
  signal N_10590 : std_logic ;
  signal N_10591 : std_logic ;
  signal N_10592 : std_logic ;
  signal N_10593 : std_logic ;
  signal N_10594 : std_logic ;
  signal N_10595 : std_logic ;
  signal N_10596 : std_logic ;
  signal N_10597 : std_logic ;
  signal N_10598 : std_logic ;
  signal N_10599 : std_logic ;
  signal N_10600 : std_logic ;
  signal N_10601 : std_logic ;
  signal N_10602 : std_logic ;
  signal N_10603 : std_logic ;
  signal N_10604 : std_logic ;
  signal N_10605 : std_logic ;
  signal N_10606 : std_logic ;
  signal N_10607 : std_logic ;
  signal N_10608 : std_logic ;
  signal N_10609 : std_logic ;
  signal N_10610 : std_logic ;
  signal N_10611 : std_logic ;
  signal N_10612 : std_logic ;
  signal N_10613 : std_logic ;
  signal N_10614 : std_logic ;
  signal N_10615 : std_logic ;
  signal N_10616 : std_logic ;
  signal N_10617 : std_logic ;
  signal N_10618 : std_logic ;
  signal N_10619 : std_logic ;
  signal N_10620 : std_logic ;
  signal N_10621 : std_logic ;
  signal N_10622 : std_logic ;
  signal N_10623 : std_logic ;
  signal N_10624 : std_logic ;
  signal N_10625 : std_logic ;
  signal N_10626 : std_logic ;
  signal N_10627 : std_logic ;
  signal N_10628 : std_logic ;
  signal N_10629 : std_logic ;
  signal N_10630 : std_logic ;
  signal N_10631 : std_logic ;
  signal R1IN_4_ADD_2_1 : std_logic ;
  signal NN_3 : std_logic ;
  signal NN_4 : std_logic ;
  signal NN_5 : std_logic ;
  signal NN_6 : std_logic ;
  signal NN_7 : std_logic ;
  signal NN_8 : std_logic ;
  signal NN_9 : std_logic ;
  signal NN_10 : std_logic ;
  signal N_10632 : std_logic ;
  signal N_10806 : std_logic ;
  signal N_10807 : std_logic ;
  signal N_10808 : std_logic ;
  signal N_10809 : std_logic ;
  signal N_10810 : std_logic ;
  signal N_10811 : std_logic ;
  signal N_10812 : std_logic ;
  signal N_10813 : std_logic ;
  signal N_10814 : std_logic ;
  signal N_10815 : std_logic ;
  signal N_10816 : std_logic ;
  signal N_10817 : std_logic ;
  signal N_10818 : std_logic ;
  signal N_10819 : std_logic ;
  signal N_10820 : std_logic ;
  signal N_10821 : std_logic ;
  signal N_10822 : std_logic ;
  signal N_10823 : std_logic ;
  signal N_10824 : std_logic ;
  signal N_10825 : std_logic ;
  signal N_10826 : std_logic ;
  signal N_10827 : std_logic ;
  signal N_10828 : std_logic ;
  signal N_10829 : std_logic ;
  signal N_10830 : std_logic ;
  signal N_10831 : std_logic ;
  signal N_10832 : std_logic ;
  signal N_10833 : std_logic ;
  signal N_10834 : std_logic ;
  signal N_10835 : std_logic ;
  signal N_10836 : std_logic ;
  signal N_10837 : std_logic ;
  signal N_10838 : std_logic ;
  signal N_10839 : std_logic ;
  signal N_10840 : std_logic ;
  signal N_10841 : std_logic ;
  signal N_10842 : std_logic ;
  signal N_10843 : std_logic ;
  signal N_10844 : std_logic ;
  signal N_10845 : std_logic ;
  signal N_10846 : std_logic ;
  signal N_10847 : std_logic ;
  signal N_10848 : std_logic ;
  signal N_1781_RETI : std_logic ;
  signal R2_PIPE_104_RET_1027 : std_logic ;
  signal N_1779_RETI : std_logic ;
  signal R2_PIPE_104_RET_1028 : std_logic ;
  signal N_1777_RETI : std_logic ;
  signal R2_PIPE_104_RET_1029 : std_logic ;
  signal N_1775_RETI : std_logic ;
  signal R2_PIPE_104_RET_1030 : std_logic ;
  signal N_1773_RETI : std_logic ;
  signal R2_PIPE_104_RET_1031 : std_logic ;
  signal N_1771_RETI : std_logic ;
  signal R2_PIPE_104_RET_1032 : std_logic ;
  signal N_1769_RETI : std_logic ;
  signal R2_PIPE_104_RET_1033 : std_logic ;
  signal N_1767_RETI : std_logic ;
  signal R2_PIPE_104_RET_1034 : std_logic ;
  signal N_1765_RETI : std_logic ;
  signal R2_PIPE_104_RET_1035 : std_logic ;
  signal N_1763_RETI : std_logic ;
  signal R2_PIPE_104_RET_1036 : std_logic ;
  signal N_1761_RETI : std_logic ;
  signal R2_PIPE_104_RET_1037 : std_logic ;
  signal N_1759_RETI : std_logic ;
  signal R2_PIPE_104_RET_1038 : std_logic ;
  signal N_1757_RETI : std_logic ;
  signal R2_PIPE_104_RET_1039 : std_logic ;
  signal N_1755_RETI : std_logic ;
  signal R2_PIPE_104_RET_1040 : std_logic ;
  signal N_1753_RETI : std_logic ;
  signal R2_PIPE_104_RET_1041 : std_logic ;
  signal N_1751_RETI : std_logic ;
  signal R2_PIPE_104_RET_1042 : std_logic ;
  signal N_1749_RETI : std_logic ;
  signal R2_PIPE_104_RET_1043 : std_logic ;
  signal N_1747_RETI : std_logic ;
  signal R2_PIPE_104_RET_1044 : std_logic ;
  signal N_1745_RETI : std_logic ;
  signal R2_PIPE_104_RET_1045 : std_logic ;
  signal N_1743_RETI : std_logic ;
  signal R2_PIPE_104_RET_1046 : std_logic ;
  signal N_1741_RETI : std_logic ;
  signal R2_PIPE_104_RET_1047 : std_logic ;
  signal N_1739_RETI : std_logic ;
  signal R2_PIPE_104_RET_1048 : std_logic ;
  signal N_1737_RETI : std_logic ;
  signal R2_PIPE_104_RET_1049 : std_logic ;
  signal N_1735_RETI : std_logic ;
  signal R2_PIPE_104_RET_1050 : std_logic ;
  signal N_1733_RETI : std_logic ;
  signal R2_PIPE_104_RET_1051 : std_logic ;
  signal N_1731_RETI : std_logic ;
  signal R2_PIPE_104_RET_1052 : std_logic ;
  signal N_1729_RETI : std_logic ;
  signal R2_PIPE_104_RET_1053 : std_logic ;
  signal N_1727_RETI : std_logic ;
  signal R2_PIPE_104_RET_1054 : std_logic ;
  signal N_1725_RETI : std_logic ;
  signal R2_PIPE_104_RET_1055 : std_logic ;
  signal N_1723_RETI : std_logic ;
  signal R2_PIPE_104_RET_1056 : std_logic ;
  signal N_1721_RETI : std_logic ;
  signal R2_PIPE_104_RET_1057 : std_logic ;
  signal N_1719_RETI : std_logic ;
  signal R2_PIPE_104_RET_1058 : std_logic ;
  signal N_1717_RETI : std_logic ;
  signal R2_PIPE_104_RET_1059 : std_logic ;
  signal N_1715_RETI : std_logic ;
  signal R2_PIPE_104_RET_1060 : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_0_RETI : std_logic ;
  signal R1IN_4_ADD_2_1_AXB_0 : std_logic ;
  signal N_10849 : std_logic ;
  signal NN_11 : std_logic ;
  component DSP48

    generic (
      AREG : integer := 0;
      BREG : integer := 0;
      CREG : integer := 0;
      PREG : integer := 0;
      MREG : integer := 0;
      SUBTRACTREG : integer := 0;
      OPMODEREG : integer := 0;
      CARRYINSELREG : integer := 0;
      CARRYINREG : integer := 0;
      B_INPUT : string := "DIRECT";
      LEGACY_MODE : string := "MULT18X18S"
    );
    port(
      A : in std_logic_vector(17 downto 0);
      B : in std_logic_vector(17 downto 0);
      C : in std_logic_vector(47 downto 0);
      BCIN : in std_logic_vector(17 downto 0);
      PCIN : in std_logic_vector(47 downto 0);
      OPMODE : in std_logic_vector(6 downto 0);
      SUBTRACT :  in std_logic;
      CARRYIN :  in std_logic;
      CARRYINSEL : in std_logic_vector(1 downto 0);
      CLK :  in std_logic;
      CEA :  in std_logic;
      CEB :  in std_logic;
      CEC :  in std_logic;
      CEP :  in std_logic;
      CEM :  in std_logic;
      CECARRYIN :  in std_logic;
      CECTRL :  in std_logic;
      CECINSUB :  in std_logic;
      RSTA :  in std_logic;
      RSTB :  in std_logic;
      RSTC :  in std_logic;
      RSTP :  in std_logic;
      RSTM :  in std_logic;
      RSTCTRL :  in std_logic;
      RSTCARRYIN :  in std_logic;
      BCOUT : out std_logic_vector(17 downto 0);
      P : out std_logic_vector(47 downto 0);
      PCOUT : out std_logic_vector(47 downto 0)  );
  end component;
begin
R1IN_ADD_2_0_AXB_1_Z5286: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(18),
  I1 => R1IN_ADD_1FF(1),
  O => R1IN_ADD_2_0_AXB_1);
R1IN_ADD_2_0_AXB_2_Z5287: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(19),
  I1 => R1IN_ADD_1FF(2),
  O => R1IN_ADD_2_0_AXB_2);
R1IN_ADD_2_0_AXB_3_Z5288: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(20),
  I1 => R1IN_ADD_1FF(3),
  O => R1IN_ADD_2_0_AXB_3);
R1IN_ADD_2_0_AXB_4_Z5289: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(21),
  I1 => R1IN_ADD_1FF(4),
  O => R1IN_ADD_2_0_AXB_4);
R1IN_ADD_2_0_AXB_5_Z5290: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(22),
  I1 => R1IN_ADD_1FF(5),
  O => R1IN_ADD_2_0_AXB_5);
R1IN_ADD_2_0_AXB_6_Z5291: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(23),
  I1 => R1IN_ADD_1FF(6),
  O => R1IN_ADD_2_0_AXB_6);
R1IN_ADD_2_0_AXB_7_Z5292: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(24),
  I1 => R1IN_ADD_1FF(7),
  O => R1IN_ADD_2_0_AXB_7);
R1IN_ADD_2_0_AXB_8_Z5293: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(25),
  I1 => R1IN_ADD_1FF(8),
  O => R1IN_ADD_2_0_AXB_8);
R1IN_ADD_2_0_AXB_9_Z5294: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(26),
  I1 => R1IN_ADD_1FF(9),
  O => R1IN_ADD_2_0_AXB_9);
R1IN_ADD_2_0_AXB_10_Z5295: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(27),
  I1 => R1IN_ADD_1FF(10),
  O => R1IN_ADD_2_0_AXB_10);
R1IN_ADD_2_0_AXB_11_Z5296: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(28),
  I1 => R1IN_ADD_1FF(11),
  O => R1IN_ADD_2_0_AXB_11);
R1IN_ADD_2_0_AXB_12_Z5297: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(29),
  I1 => R1IN_ADD_1FF(12),
  O => R1IN_ADD_2_0_AXB_12);
R1IN_ADD_2_0_AXB_13_Z5298: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(30),
  I1 => R1IN_ADD_1FF(13),
  O => R1IN_ADD_2_0_AXB_13);
R1IN_ADD_2_0_AXB_14_Z5299: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(31),
  I1 => R1IN_ADD_1FF(14),
  O => R1IN_ADD_2_0_AXB_14);
R1IN_ADD_2_0_AXB_15_Z5300: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(32),
  I1 => R1IN_ADD_1FF(15),
  O => R1IN_ADD_2_0_AXB_15);
R1IN_ADD_2_0_AXB_16_Z5301: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_1FF(33),
  I1 => R1IN_ADD_1FF(16),
  O => R1IN_ADD_2_0_AXB_16);
R1IN_ADD_2_0_AXB_17_Z5302: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(0),
  I1 => R1IN_ADD_1FF(17),
  O => R1IN_ADD_2_0_AXB_17);
R1IN_ADD_2_0_AXB_18_Z5303: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(1),
  I1 => R1IN_ADD_1FF(18),
  O => R1IN_ADD_2_0_AXB_18);
R1IN_ADD_2_0_AXB_19_Z5304: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(2),
  I1 => R1IN_ADD_1FF(19),
  O => R1IN_ADD_2_0_AXB_19);
R1IN_ADD_2_0_AXB_20_Z5305: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(3),
  I1 => R1IN_ADD_1FF(20),
  O => R1IN_ADD_2_0_AXB_20);
R1IN_ADD_2_0_AXB_21_Z5306: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(4),
  I1 => R1IN_ADD_1FF(21),
  O => R1IN_ADD_2_0_AXB_21);
R1IN_ADD_2_0_AXB_22_Z5307: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(5),
  I1 => R1IN_ADD_1FF(22),
  O => R1IN_ADD_2_0_AXB_22);
R1IN_ADD_2_0_AXB_23_Z5308: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(6),
  I1 => R1IN_ADD_1FF(23),
  O => R1IN_ADD_2_0_AXB_23);
R1IN_ADD_2_0_AXB_24_Z5309: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(7),
  I1 => R1IN_ADD_1FF(24),
  O => R1IN_ADD_2_0_AXB_24);
R1IN_ADD_2_0_AXB_25_Z5310: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(8),
  I1 => R1IN_ADD_1FF(25),
  O => R1IN_ADD_2_0_AXB_25);
R1IN_ADD_2_0_AXB_26_Z5311: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(9),
  I1 => R1IN_ADD_1FF(26),
  O => R1IN_ADD_2_0_AXB_26);
R1IN_ADD_2_0_AXB_27_Z5312: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(10),
  I1 => R1IN_ADD_1FF(27),
  O => R1IN_ADD_2_0_AXB_27);
R1IN_ADD_2_0_AXB_28_Z5313: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(11),
  I1 => R1IN_ADD_1FF(28),
  O => R1IN_ADD_2_0_AXB_28);
R1IN_ADD_2_0_AXB_29_Z5314: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(12),
  I1 => R1IN_ADD_1FF(29),
  O => R1IN_ADD_2_0_AXB_29);
R1IN_ADD_2_0_AXB_30_Z5315: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(13),
  I1 => R1IN_ADD_1FF(30),
  O => R1IN_ADD_2_0_AXB_30);
R1IN_ADD_2_0_AXB_31_Z5316: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(14),
  I1 => R1IN_ADD_1FF(31),
  O => R1IN_ADD_2_0_AXB_31);
R1IN_ADD_2_0_AXB_32_Z5317: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4FF(15),
  I1 => R1IN_ADD_1FF(32),
  O => R1IN_ADD_2_0_AXB_32);
R1IN_ADD_2_0_AXB_33_Z5318: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4FF(16),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_18,
  I2 => R2_PIPE_138_RET,
  I3 => R2_PIPE_138_RET_1,
  O => R1IN_ADD_2_0_AXB_33);
R1IN_ADD_2_0_AXB_34_Z5319: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(17),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_17,
  I2 => R2_PIPE_139_RET,
  I3 => R2_PIPE_139_RET_1,
  O => R1IN_ADD_2_0_AXB_34);
R1IN_ADD_2_0_AXB_35_Z5320: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(18),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_16,
  I2 => R2_PIPE_140_RET,
  I3 => R2_PIPE_140_RET_1,
  O => R1IN_ADD_2_0_AXB_35);
R1IN_ADD_2_0_AXB_36_Z5321: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(19),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_15,
  I2 => R2_PIPE_141_RET,
  I3 => R2_PIPE_141_RET_1,
  O => R1IN_ADD_2_0_AXB_36);
R1IN_ADD_2_0_AXB_37_Z5322: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(20),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_14,
  I2 => R2_PIPE_142_RET,
  I3 => R2_PIPE_142_RET_1,
  O => R1IN_ADD_2_0_AXB_37);
R1IN_ADD_2_0_AXB_38_Z5323: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(21),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_13,
  I2 => R2_PIPE_143_RET,
  I3 => R2_PIPE_143_RET_1,
  O => R1IN_ADD_2_0_AXB_38);
R1IN_ADD_2_0_AXB_39_Z5324: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(22),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_12,
  I2 => R2_PIPE_144_RET,
  I3 => R2_PIPE_144_RET_1,
  O => R1IN_ADD_2_0_AXB_39);
R1IN_ADD_2_0_AXB_40_Z5325: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(23),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_11,
  I2 => R2_PIPE_145_RET,
  I3 => R2_PIPE_145_RET_1,
  O => R1IN_ADD_2_0_AXB_40);
R1IN_ADD_2_0_AXB_41_Z5326: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(24),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_10,
  I2 => R2_PIPE_146_RET,
  I3 => R2_PIPE_146_RET_1,
  O => R1IN_ADD_2_0_AXB_41);
R1IN_ADD_2_0_AXB_42_Z5327: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(25),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_9,
  I2 => R2_PIPE_147_RET,
  I3 => R2_PIPE_147_RET_1,
  O => R1IN_ADD_2_0_AXB_42);
R1IN_ADD_2_0_AXB_43_Z5328: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(26),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_8,
  I2 => R2_PIPE_148_RET,
  I3 => R2_PIPE_148_RET_1,
  O => R1IN_ADD_2_0_AXB_43);
R1IN_ADD_2_0_AXB_44_Z5329: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(27),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_7,
  I2 => R2_PIPE_149_RET,
  I3 => R2_PIPE_149_RET_1,
  O => R1IN_ADD_2_0_AXB_44);
R1IN_ADD_2_0_AXB_45_Z5330: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(28),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_6,
  I2 => R2_PIPE_150_RET,
  I3 => R2_PIPE_150_RET_1,
  O => R1IN_ADD_2_0_AXB_45);
R1IN_ADD_2_0_AXB_46_Z5331: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(29),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_5,
  I2 => R2_PIPE_151_RET,
  I3 => R2_PIPE_151_RET_1,
  O => R1IN_ADD_2_0_AXB_46);
R1IN_ADD_2_0_AXB_47_Z5332: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(30),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_4,
  I2 => R2_PIPE_152_RET,
  I3 => R2_PIPE_152_RET_1,
  O => R1IN_ADD_2_0_AXB_47);
R1IN_ADD_2_0_AXB_48_Z5333: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(31),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_3,
  I2 => R2_PIPE_153_RET,
  I3 => R2_PIPE_153_RET_1,
  O => R1IN_ADD_2_0_AXB_48);
R1IN_ADD_2_0_AXB_49_Z5334: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(32),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_2,
  I2 => R2_PIPE_154_RET,
  I3 => R2_PIPE_154_RET_1,
  O => R1IN_ADD_2_0_AXB_49);
R1IN_ADD_2_0_AXB_50_Z5335: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(33),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_1,
  I2 => R2_PIPE_155_RET,
  I3 => R2_PIPE_155_RET_1,
  O => R1IN_ADD_2_0_AXB_50);
R1IN_ADD_2_0_AXB_51_Z5336: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(34),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_0,
  I2 => R2_PIPE_156_RET,
  I3 => R2_PIPE_156_RET_1,
  O => R1IN_ADD_2_0_AXB_51);
R1IN_ADD_2_0_AXB_52_Z5337: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(35),
  I1 => R1IN_ADD_1_0_CRY_31_RETO,
  I2 => R2_PIPE_157_RET,
  I3 => R2_PIPE_157_RET_1,
  O => R1IN_ADD_2_0_AXB_52);
R1IN_ADD_2_1_AXB_1_Z5338: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(37),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_25,
  I2 => R2_PIPE_159_RET,
  I3 => R2_PIPE_159_RET_1,
  O => R1IN_ADD_2_1_AXB_1);
R1IN_ADD_2_1_AXB_2_Z5339: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(38),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_24,
  I2 => R2_PIPE_160_RET,
  I3 => R2_PIPE_160_RET_1,
  O => R1IN_ADD_2_1_AXB_2);
R1IN_ADD_2_1_AXB_3_Z5340: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(39),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_23,
  I2 => R2_PIPE_161_RET,
  I3 => R2_PIPE_161_RET_1,
  O => R1IN_ADD_2_1_AXB_3);
R1IN_ADD_2_1_AXB_4_Z5341: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(40),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_22,
  I2 => R2_PIPE_162_RET,
  I3 => R2_PIPE_162_RET_1,
  O => R1IN_ADD_2_1_AXB_4);
R1IN_ADD_2_1_AXB_5_Z5342: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(41),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_21,
  I2 => R2_PIPE_163_RET,
  I3 => R2_PIPE_163_RET_1,
  O => R1IN_ADD_2_1_AXB_5);
R1IN_ADD_2_1_AXB_6_Z5343: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(42),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_20,
  I2 => R2_PIPE_164_RET,
  I3 => R2_PIPE_164_RET_1,
  O => R1IN_ADD_2_1_AXB_6);
R1IN_ADD_2_1_AXB_7_Z5344: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(43),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_19,
  I2 => R2_PIPE_165_RET,
  I3 => R2_PIPE_165_RET_1,
  O => R1IN_ADD_2_1_AXB_7);
R1IN_ADD_2_1_AXB_8_Z5345: LUT4 
generic map(
  INIT => X"596A"
)
port map (
  I0 => R1IN_4F(44),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_27,
  I2 => R1IN_ADD_1_1_0_CRY_28_RETO,
  I3 => R1IN_ADD_1_1_CRY_28_RETO,
  O => R1IN_ADD_2_1_AXB_8);
R1IN_ADD_2_1_AXB_9_Z5346: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4F(45),
  O => R1IN_ADD_2_1_AXB_9);
R1IN_ADD_2_1_AXB_10_Z5347: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4F(46),
  O => R1IN_ADD_2_1_AXB_10);
R1IN_ADD_2_1_AXB_11_Z5348: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4F(47),
  O => R1IN_ADD_2_1_AXB_11);
R1IN_ADD_2_1_AXB_12_Z5349: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4F(48),
  O => R1IN_ADD_2_1_AXB_12);
R1IN_ADD_2_1_AXB_13_Z5350: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4F(49),
  O => R1IN_ADD_2_1_AXB_13);
R1IN_ADD_2_1_AXB_14_Z5351: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4F(50),
  O => R1IN_ADD_2_1_AXB_14);
R1IN_ADD_2_1_AXB_15_Z5352: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4F(51),
  O => R1IN_ADD_2_1_AXB_15);
R1IN_ADD_2_1_AXB_16_Z5353: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4F(52),
  O => R1IN_ADD_2_1_AXB_16);
R1IN_ADD_2_1_AXB_17_Z5354: LUT3 
generic map(
  INIT => X"72"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_32,
  I1 => R1IN_4_ADD_2_1_0_AXB_0_RETO,
  I2 => R1IN_4_ADD_2_1_AXB_0,
  O => R1IN_ADD_2_1_AXB_17);
R1IN_ADD_2_1_AXB_18_Z5355: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4(54),
  O => R1IN_ADD_2_1_AXB_18);
R1IN_ADD_2_1_AXB_19_Z5356: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_31,
  I1 => R2_PIPE_104_RET_123,
  I2 => R2_PIPE_104_RET_1059,
  O => R1IN_ADD_2_1_AXB_19);
R1IN_ADD_2_1_AXB_20_Z5357: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_30,
  I1 => R2_PIPE_104_RET_122,
  I2 => R2_PIPE_104_RET_1058,
  O => R1IN_ADD_2_1_AXB_20);
R1IN_ADD_2_1_AXB_21_Z5358: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_29,
  I1 => R2_PIPE_104_RET_121,
  I2 => R2_PIPE_104_RET_1057,
  O => R1IN_ADD_2_1_AXB_21);
R1IN_ADD_2_1_AXB_22_Z5359: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_28,
  I1 => R2_PIPE_104_RET_120,
  I2 => R2_PIPE_104_RET_1056,
  O => R1IN_ADD_2_1_AXB_22);
R1IN_ADD_2_1_AXB_23_Z5360: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_27,
  I1 => R2_PIPE_104_RET_119,
  I2 => R2_PIPE_104_RET_1055,
  O => R1IN_ADD_2_1_AXB_23);
R1IN_ADD_2_1_AXB_24_Z5361: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_26,
  I1 => R2_PIPE_104_RET_118,
  I2 => R2_PIPE_104_RET_1054,
  O => R1IN_ADD_2_1_AXB_24);
R1IN_ADD_2_1_AXB_25_Z5362: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_25,
  I1 => R2_PIPE_104_RET_117,
  I2 => R2_PIPE_104_RET_1053,
  O => R1IN_ADD_2_1_AXB_25);
R1IN_ADD_2_1_AXB_26_Z5363: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_24,
  I1 => R2_PIPE_104_RET_116,
  I2 => R2_PIPE_104_RET_1052,
  O => R1IN_ADD_2_1_AXB_26);
R1IN_ADD_2_1_AXB_27_Z5364: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_23,
  I1 => R2_PIPE_104_RET_115,
  I2 => R2_PIPE_104_RET_1051,
  O => R1IN_ADD_2_1_AXB_27);
R1IN_ADD_2_1_AXB_28_Z5365: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_22,
  I1 => R2_PIPE_104_RET_114,
  I2 => R2_PIPE_104_RET_1050,
  O => R1IN_ADD_2_1_AXB_28);
R1IN_ADD_2_1_AXB_29_Z5366: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_21,
  I1 => R2_PIPE_104_RET_113,
  I2 => R2_PIPE_104_RET_1049,
  O => R1IN_ADD_2_1_AXB_29);
R1IN_ADD_2_1_AXB_30_Z5367: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_20,
  I1 => R2_PIPE_104_RET_112,
  I2 => R2_PIPE_104_RET_1048,
  O => R1IN_ADD_2_1_AXB_30);
R1IN_ADD_2_1_AXB_31_Z5368: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_19,
  I1 => R2_PIPE_104_RET_111,
  I2 => R2_PIPE_104_RET_1047,
  O => R1IN_ADD_2_1_AXB_31);
R1IN_ADD_2_1_AXB_32_Z5369: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_18,
  I1 => R2_PIPE_104_RET_110,
  I2 => R2_PIPE_104_RET_1046,
  O => R1IN_ADD_2_1_AXB_32);
R1IN_ADD_2_1_AXB_33_Z5370: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_17,
  I1 => R2_PIPE_104_RET_109,
  I2 => R2_PIPE_104_RET_1045,
  O => R1IN_ADD_2_1_AXB_33);
R1IN_ADD_2_1_AXB_34_Z5371: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_16,
  I1 => R2_PIPE_104_RET_108,
  I2 => R2_PIPE_104_RET_1044,
  O => R1IN_ADD_2_1_AXB_34);
R1IN_ADD_2_1_AXB_35_Z5372: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_15,
  I1 => R2_PIPE_104_RET_107,
  I2 => R2_PIPE_104_RET_1043,
  O => R1IN_ADD_2_1_AXB_35);
R1IN_ADD_2_1_AXB_36_Z5373: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_14,
  I1 => R2_PIPE_104_RET_106,
  I2 => R2_PIPE_104_RET_1042,
  O => R1IN_ADD_2_1_AXB_36);
R1IN_ADD_2_1_AXB_37_Z5374: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_13,
  I1 => R2_PIPE_104_RET_105,
  I2 => R2_PIPE_104_RET_1041,
  O => R1IN_ADD_2_1_AXB_37);
R1IN_ADD_2_1_AXB_38_Z5375: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_12,
  I1 => R2_PIPE_104_RET_104,
  I2 => R2_PIPE_104_RET_1040,
  O => R1IN_ADD_2_1_AXB_38);
R1IN_ADD_2_1_AXB_39_Z5376: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_11,
  I1 => R2_PIPE_104_RET_103,
  I2 => R2_PIPE_104_RET_1039,
  O => R1IN_ADD_2_1_AXB_39);
R1IN_ADD_2_1_AXB_40_Z5377: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_10,
  I1 => R2_PIPE_104_RET_102,
  I2 => R2_PIPE_104_RET_1038,
  O => R1IN_ADD_2_1_AXB_40);
R1IN_ADD_2_1_AXB_41_Z5378: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_9,
  I1 => R2_PIPE_104_RET_101,
  I2 => R2_PIPE_104_RET_1037,
  O => R1IN_ADD_2_1_AXB_41);
R1IN_ADD_2_1_AXB_42_Z5379: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_8,
  I1 => R2_PIPE_104_RET_100,
  I2 => R2_PIPE_104_RET_1036,
  O => R1IN_ADD_2_1_AXB_42);
R1IN_ADD_2_1_AXB_43_Z5380: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_7,
  I1 => R2_PIPE_104_RET_99,
  I2 => R2_PIPE_104_RET_1035,
  O => R1IN_ADD_2_1_AXB_43);
R1IN_ADD_2_1_AXB_44_Z5381: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_6,
  I1 => R2_PIPE_104_RET_98,
  I2 => R2_PIPE_104_RET_1034,
  O => R1IN_ADD_2_1_AXB_44);
R1IN_ADD_2_1_AXB_45_Z5382: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_5,
  I1 => R2_PIPE_104_RET_97,
  I2 => R2_PIPE_104_RET_1033,
  O => R1IN_ADD_2_1_AXB_45);
R1IN_ADD_2_1_AXB_46_Z5383: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_4,
  I1 => R2_PIPE_104_RET_96,
  I2 => R2_PIPE_104_RET_1032,
  O => R1IN_ADD_2_1_AXB_46);
R1IN_ADD_2_1_AXB_47_Z5384: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_3,
  I1 => R2_PIPE_104_RET_95,
  I2 => R2_PIPE_104_RET_1031,
  O => R1IN_ADD_2_1_AXB_47);
R1IN_ADD_2_1_AXB_48_Z5385: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_2,
  I1 => R2_PIPE_104_RET_94,
  I2 => R2_PIPE_104_RET_1030,
  O => R1IN_ADD_2_1_AXB_48);
R1IN_ADD_2_1_AXB_49_Z5386: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_1,
  I1 => R2_PIPE_104_RET_93,
  I2 => R2_PIPE_104_RET_1029,
  O => R1IN_ADD_2_1_AXB_49);
R1IN_ADD_2_1_AXB_50_Z5387: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_0,
  I1 => R2_PIPE_104_RET_49,
  I2 => R2_PIPE_104_RET_1028,
  O => R1IN_ADD_2_1_AXB_50);
R1IN_ADD_2_1_0_AXB_1_Z5388: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(37),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_25,
  I2 => R2_PIPE_159_RET,
  I3 => R2_PIPE_159_RET_1,
  O => R1IN_ADD_2_1_0_AXB_1);
R1IN_ADD_2_1_0_AXB_2_Z5389: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(38),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_24,
  I2 => R2_PIPE_160_RET,
  I3 => R2_PIPE_160_RET_1,
  O => R1IN_ADD_2_1_0_AXB_2);
R1IN_ADD_2_1_0_AXB_3_Z5390: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(39),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_23,
  I2 => R2_PIPE_161_RET,
  I3 => R2_PIPE_161_RET_1,
  O => R1IN_ADD_2_1_0_AXB_3);
R1IN_ADD_2_1_0_AXB_4_Z5391: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(40),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_22,
  I2 => R2_PIPE_162_RET,
  I3 => R2_PIPE_162_RET_1,
  O => R1IN_ADD_2_1_0_AXB_4);
R1IN_ADD_2_1_0_AXB_5_Z5392: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(41),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_21,
  I2 => R2_PIPE_163_RET,
  I3 => R2_PIPE_163_RET_1,
  O => R1IN_ADD_2_1_0_AXB_5);
R1IN_ADD_2_1_0_AXB_6_Z5393: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(42),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_20,
  I2 => R2_PIPE_164_RET,
  I3 => R2_PIPE_164_RET_1,
  O => R1IN_ADD_2_1_0_AXB_6);
R1IN_ADD_2_1_0_AXB_7_Z5394: LUT4 
generic map(
  INIT => X"569A"
)
port map (
  I0 => R1IN_4F(43),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_19,
  I2 => R2_PIPE_165_RET,
  I3 => R2_PIPE_165_RET_1,
  O => R1IN_ADD_2_1_0_AXB_7);
R1IN_ADD_2_1_0_AXB_8_Z5395: LUT4 
generic map(
  INIT => X"596A"
)
port map (
  I0 => R1IN_4F(44),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_27,
  I2 => R1IN_ADD_1_1_0_CRY_28_RETO,
  I3 => R1IN_ADD_1_1_CRY_28_RETO,
  O => R1IN_ADD_2_1_0_AXB_8);
R1IN_ADD_2_1_0_AXB_9_Z5396: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4F(45),
  O => R1IN_ADD_2_1_0_AXB_9);
R1IN_ADD_2_1_0_AXB_10_Z5397: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4F(46),
  O => R1IN_ADD_2_1_0_AXB_10);
R1IN_ADD_2_1_0_AXB_11_Z5398: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4F(47),
  O => R1IN_ADD_2_1_0_AXB_11);
R1IN_ADD_2_1_0_AXB_12_Z5399: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4F(48),
  O => R1IN_ADD_2_1_0_AXB_12);
R1IN_ADD_2_1_0_AXB_13_Z5400: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4F(49),
  O => R1IN_ADD_2_1_0_AXB_13);
R1IN_ADD_2_1_0_AXB_14_Z5401: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4F(50),
  O => R1IN_ADD_2_1_0_AXB_14);
R1IN_ADD_2_1_0_AXB_15_Z5402: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4F(51),
  O => R1IN_ADD_2_1_0_AXB_15);
R1IN_ADD_2_1_0_AXB_16_Z5403: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4F(52),
  O => R1IN_ADD_2_1_0_AXB_16);
R1IN_ADD_2_1_0_AXB_17_Z5404: LUT3 
generic map(
  INIT => X"72"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_32,
  I1 => R1IN_4_ADD_2_1_0_AXB_0_RETO,
  I2 => R1IN_4_ADD_2_1_AXB_0,
  O => R1IN_ADD_2_1_0_AXB_17);
R1IN_ADD_2_1_0_AXB_18_Z5405: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4(54),
  O => R1IN_ADD_2_1_0_AXB_18);
R1IN_ADD_2_1_0_AXB_19_Z5406: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_31,
  I1 => R2_PIPE_104_RET_123,
  I2 => R2_PIPE_104_RET_1059,
  O => R1IN_ADD_2_1_0_AXB_19);
R1IN_ADD_2_1_0_AXB_20_Z5407: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_30,
  I1 => R2_PIPE_104_RET_122,
  I2 => R2_PIPE_104_RET_1058,
  O => R1IN_ADD_2_1_0_AXB_20);
R1IN_ADD_2_1_0_AXB_21_Z5408: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_29,
  I1 => R2_PIPE_104_RET_121,
  I2 => R2_PIPE_104_RET_1057,
  O => R1IN_ADD_2_1_0_AXB_21);
R1IN_ADD_2_1_0_AXB_22_Z5409: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_28,
  I1 => R2_PIPE_104_RET_120,
  I2 => R2_PIPE_104_RET_1056,
  O => R1IN_ADD_2_1_0_AXB_22);
R1IN_ADD_2_1_0_AXB_23_Z5410: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_27,
  I1 => R2_PIPE_104_RET_119,
  I2 => R2_PIPE_104_RET_1055,
  O => R1IN_ADD_2_1_0_AXB_23);
R1IN_ADD_2_1_0_AXB_24_Z5411: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_26,
  I1 => R2_PIPE_104_RET_118,
  I2 => R2_PIPE_104_RET_1054,
  O => R1IN_ADD_2_1_0_AXB_24);
R1IN_ADD_2_1_0_AXB_25_Z5412: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_25,
  I1 => R2_PIPE_104_RET_117,
  I2 => R2_PIPE_104_RET_1053,
  O => R1IN_ADD_2_1_0_AXB_25);
R1IN_ADD_2_1_0_AXB_26_Z5413: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_24,
  I1 => R2_PIPE_104_RET_116,
  I2 => R2_PIPE_104_RET_1052,
  O => R1IN_ADD_2_1_0_AXB_26);
R1IN_ADD_2_1_0_AXB_27_Z5414: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_23,
  I1 => R2_PIPE_104_RET_115,
  I2 => R2_PIPE_104_RET_1051,
  O => R1IN_ADD_2_1_0_AXB_27);
R1IN_ADD_2_1_0_AXB_28_Z5415: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_22,
  I1 => R2_PIPE_104_RET_114,
  I2 => R2_PIPE_104_RET_1050,
  O => R1IN_ADD_2_1_0_AXB_28);
R1IN_ADD_2_1_0_AXB_29_Z5416: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_21,
  I1 => R2_PIPE_104_RET_113,
  I2 => R2_PIPE_104_RET_1049,
  O => R1IN_ADD_2_1_0_AXB_29);
R1IN_ADD_2_1_0_AXB_30_Z5417: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_20,
  I1 => R2_PIPE_104_RET_112,
  I2 => R2_PIPE_104_RET_1048,
  O => R1IN_ADD_2_1_0_AXB_30);
R1IN_ADD_2_1_0_AXB_31_Z5418: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_19,
  I1 => R2_PIPE_104_RET_111,
  I2 => R2_PIPE_104_RET_1047,
  O => R1IN_ADD_2_1_0_AXB_31);
R1IN_ADD_2_1_0_AXB_32_Z5419: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_18,
  I1 => R2_PIPE_104_RET_110,
  I2 => R2_PIPE_104_RET_1046,
  O => R1IN_ADD_2_1_0_AXB_32);
R1IN_ADD_2_1_0_AXB_33_Z5420: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_17,
  I1 => R2_PIPE_104_RET_109,
  I2 => R2_PIPE_104_RET_1045,
  O => R1IN_ADD_2_1_0_AXB_33);
R1IN_ADD_2_1_0_AXB_34_Z5421: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_16,
  I1 => R2_PIPE_104_RET_108,
  I2 => R2_PIPE_104_RET_1044,
  O => R1IN_ADD_2_1_0_AXB_34);
R1IN_ADD_2_1_0_AXB_35_Z5422: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_15,
  I1 => R2_PIPE_104_RET_107,
  I2 => R2_PIPE_104_RET_1043,
  O => R1IN_ADD_2_1_0_AXB_35);
R1IN_ADD_2_1_0_AXB_36_Z5423: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_14,
  I1 => R2_PIPE_104_RET_106,
  I2 => R2_PIPE_104_RET_1042,
  O => R1IN_ADD_2_1_0_AXB_36);
R1IN_ADD_2_1_0_AXB_37_Z5424: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_13,
  I1 => R2_PIPE_104_RET_105,
  I2 => R2_PIPE_104_RET_1041,
  O => R1IN_ADD_2_1_0_AXB_37);
R1IN_ADD_2_1_0_AXB_38_Z5425: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_12,
  I1 => R2_PIPE_104_RET_104,
  I2 => R2_PIPE_104_RET_1040,
  O => R1IN_ADD_2_1_0_AXB_38);
R1IN_ADD_2_1_0_AXB_39_Z5426: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_11,
  I1 => R2_PIPE_104_RET_103,
  I2 => R2_PIPE_104_RET_1039,
  O => R1IN_ADD_2_1_0_AXB_39);
R1IN_ADD_2_1_0_AXB_40_Z5427: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_10,
  I1 => R2_PIPE_104_RET_102,
  I2 => R2_PIPE_104_RET_1038,
  O => R1IN_ADD_2_1_0_AXB_40);
R1IN_ADD_2_1_0_AXB_41_Z5428: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_9,
  I1 => R2_PIPE_104_RET_101,
  I2 => R2_PIPE_104_RET_1037,
  O => R1IN_ADD_2_1_0_AXB_41);
R1IN_ADD_2_1_0_AXB_42_Z5429: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_8,
  I1 => R2_PIPE_104_RET_100,
  I2 => R2_PIPE_104_RET_1036,
  O => R1IN_ADD_2_1_0_AXB_42);
R1IN_ADD_2_1_0_AXB_43_Z5430: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_7,
  I1 => R2_PIPE_104_RET_99,
  I2 => R2_PIPE_104_RET_1035,
  O => R1IN_ADD_2_1_0_AXB_43);
R1IN_ADD_2_1_0_AXB_44_Z5431: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_6,
  I1 => R2_PIPE_104_RET_98,
  I2 => R2_PIPE_104_RET_1034,
  O => R1IN_ADD_2_1_0_AXB_44);
R1IN_ADD_2_1_0_AXB_45_Z5432: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_5,
  I1 => R2_PIPE_104_RET_97,
  I2 => R2_PIPE_104_RET_1033,
  O => R1IN_ADD_2_1_0_AXB_45);
R1IN_ADD_2_1_0_AXB_46_Z5433: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_4,
  I1 => R2_PIPE_104_RET_96,
  I2 => R2_PIPE_104_RET_1032,
  O => R1IN_ADD_2_1_0_AXB_46);
R1IN_ADD_2_1_0_AXB_47_Z5434: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_3,
  I1 => R2_PIPE_104_RET_95,
  I2 => R2_PIPE_104_RET_1031,
  O => R1IN_ADD_2_1_0_AXB_47);
R1IN_ADD_2_1_0_AXB_48_Z5435: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_2,
  I1 => R2_PIPE_104_RET_94,
  I2 => R2_PIPE_104_RET_1030,
  O => R1IN_ADD_2_1_0_AXB_48);
R1IN_ADD_2_1_0_AXB_49_Z5436: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_1,
  I1 => R2_PIPE_104_RET_93,
  I2 => R2_PIPE_104_RET_1029,
  O => R1IN_ADD_2_1_0_AXB_49);
R1IN_ADD_2_1_0_AXB_50_Z5437: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO_0,
  I1 => R2_PIPE_104_RET_49,
  I2 => R2_PIPE_104_RET_1028,
  O => R1IN_ADD_2_1_0_AXB_50);
R1IN_3_ADD_1_AXB_1_Z5438: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F(18),
  I1 => R1IN_3_2F(1),
  O => R1IN_3_ADD_1_AXB_1);
R1IN_3_ADD_1_AXB_2_Z5439: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F(19),
  I1 => R1IN_3_2F(2),
  O => R1IN_3_ADD_1_AXB_2);
R1IN_3_ADD_1_AXB_3_Z5440: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F(20),
  I1 => R1IN_3_2F(3),
  O => R1IN_3_ADD_1_AXB_3);
R1IN_3_ADD_1_AXB_4_Z5441: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F(21),
  I1 => R1IN_3_2F(4),
  O => R1IN_3_ADD_1_AXB_4);
R1IN_3_ADD_1_AXB_5_Z5442: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F(22),
  I1 => R1IN_3_2F(5),
  O => R1IN_3_ADD_1_AXB_5);
R1IN_3_ADD_1_AXB_6_Z5443: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F(23),
  I1 => R1IN_3_2F(6),
  O => R1IN_3_ADD_1_AXB_6);
R1IN_3_ADD_1_AXB_7_Z5444: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F(24),
  I1 => R1IN_3_2F(7),
  O => R1IN_3_ADD_1_AXB_7);
R1IN_3_ADD_1_AXB_8_Z5445: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F(25),
  I1 => R1IN_3_2F(8),
  O => R1IN_3_ADD_1_AXB_8);
R1IN_3_ADD_1_AXB_9_Z5446: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F(26),
  I1 => R1IN_3_2F(9),
  O => R1IN_3_ADD_1_AXB_9);
R1IN_3_ADD_1_AXB_10_Z5447: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F(27),
  I1 => R1IN_3_2F(10),
  O => R1IN_3_ADD_1_AXB_10);
R1IN_3_ADD_1_AXB_11_Z5448: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F(28),
  I1 => R1IN_3_2F(11),
  O => R1IN_3_ADD_1_AXB_11);
R1IN_3_ADD_1_AXB_12_Z5449: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F(29),
  I1 => R1IN_3_2F(12),
  O => R1IN_3_ADD_1_AXB_12);
R1IN_3_ADD_1_AXB_13_Z5450: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F(30),
  I1 => R1IN_3_2F(13),
  O => R1IN_3_ADD_1_AXB_13);
R1IN_3_ADD_1_AXB_14_Z5451: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F(31),
  I1 => R1IN_3_2F(14),
  O => R1IN_3_ADD_1_AXB_14);
R1IN_3_ADD_1_AXB_15_Z5452: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F(32),
  I1 => R1IN_3_2F(15),
  O => R1IN_3_ADD_1_AXB_15);
R1IN_3_ADD_1_AXB_16_Z5453: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F(33),
  I1 => R1IN_3_2F(16),
  O => R1IN_3_ADD_1_AXB_16);
R1IN_3_ADD_1_AXB_17_Z5454: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(17),
  O => R1IN_3_ADD_1_AXB_17);
R1IN_3_ADD_1_AXB_18_Z5455: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(18),
  O => R1IN_3_ADD_1_AXB_18);
R1IN_3_ADD_1_AXB_19_Z5456: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(19),
  O => R1IN_3_ADD_1_AXB_19);
R1IN_3_ADD_1_AXB_20_Z5457: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(20),
  O => R1IN_3_ADD_1_AXB_20);
R1IN_3_ADD_1_AXB_21_Z5458: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(21),
  O => R1IN_3_ADD_1_AXB_21);
R1IN_3_ADD_1_AXB_22_Z5459: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(22),
  O => R1IN_3_ADD_1_AXB_22);
R1IN_3_ADD_1_AXB_23_Z5460: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(23),
  O => R1IN_3_ADD_1_AXB_23);
R1IN_3_ADD_1_AXB_24_Z5461: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(24),
  O => R1IN_3_ADD_1_AXB_24);
R1IN_3_ADD_1_AXB_25_Z5462: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(25),
  O => R1IN_3_ADD_1_AXB_25);
R1IN_3_ADD_1_AXB_26_Z5463: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(26),
  O => R1IN_3_ADD_1_AXB_26);
R1IN_3_ADD_1_AXB_27_Z5464: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(27),
  O => R1IN_3_ADD_1_AXB_27);
R1IN_3_ADD_1_AXB_28_Z5465: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(28),
  O => R1IN_3_ADD_1_AXB_28);
R1IN_3_ADD_1_AXB_29_Z5466: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(29),
  O => R1IN_3_ADD_1_AXB_29);
R1IN_3_ADD_1_AXB_30_Z5467: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(30),
  O => R1IN_3_ADD_1_AXB_30);
R1IN_3_ADD_1_AXB_31_Z5468: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(31),
  O => R1IN_3_ADD_1_AXB_31);
R1IN_3_ADD_1_AXB_32_Z5469: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(32),
  O => R1IN_3_ADD_1_AXB_32);
R1IN_3_ADD_1_AXB_33_Z5470: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(33),
  O => R1IN_3_ADD_1_AXB_33);
R1IN_3_ADD_1_AXB_34_Z5471: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(34),
  O => R1IN_3_ADD_1_AXB_34);
R1IN_3_ADD_1_AXB_35_Z5472: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(35),
  O => R1IN_3_ADD_1_AXB_35);
R1IN_3_ADD_1_AXB_36_Z5473: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(36),
  O => R1IN_3_ADD_1_AXB_36);
R1IN_3_ADD_1_AXB_37_Z5474: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(37),
  O => R1IN_3_ADD_1_AXB_37);
R1IN_3_ADD_1_AXB_38_Z5475: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(38),
  O => R1IN_3_ADD_1_AXB_38);
R1IN_3_ADD_1_AXB_39_Z5476: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(39),
  O => R1IN_3_ADD_1_AXB_39);
R1IN_3_ADD_1_AXB_40_Z5477: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(40),
  O => R1IN_3_ADD_1_AXB_40);
R1IN_3_ADD_1_AXB_41_Z5478: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(41),
  O => R1IN_3_ADD_1_AXB_41);
R1IN_3_ADD_1_AXB_42_Z5479: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(42),
  O => R1IN_3_ADD_1_AXB_42);
R1IN_2_ADD_1_AXB_0: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F(17),
  I1 => R1IN_2_ADD_1,
  O => R1IN_2(17));
R1IN_2_ADD_1_AXB_1_Z5481: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F(18),
  I1 => R1IN_2_2F(1),
  O => R1IN_2_ADD_1_AXB_1);
R1IN_2_ADD_1_AXB_2_Z5482: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F(19),
  I1 => R1IN_2_2F(2),
  O => R1IN_2_ADD_1_AXB_2);
R1IN_2_ADD_1_AXB_3_Z5483: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F(20),
  I1 => R1IN_2_2F(3),
  O => R1IN_2_ADD_1_AXB_3);
R1IN_2_ADD_1_AXB_4_Z5484: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F(21),
  I1 => R1IN_2_2F(4),
  O => R1IN_2_ADD_1_AXB_4);
R1IN_2_ADD_1_AXB_5_Z5485: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F(22),
  I1 => R1IN_2_2F(5),
  O => R1IN_2_ADD_1_AXB_5);
R1IN_2_ADD_1_AXB_6_Z5486: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F(23),
  I1 => R1IN_2_2F(6),
  O => R1IN_2_ADD_1_AXB_6);
R1IN_2_ADD_1_AXB_7_Z5487: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F(24),
  I1 => R1IN_2_2F(7),
  O => R1IN_2_ADD_1_AXB_7);
R1IN_2_ADD_1_AXB_8_Z5488: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F(25),
  I1 => R1IN_2_2F(8),
  O => R1IN_2_ADD_1_AXB_8);
R1IN_2_ADD_1_AXB_9_Z5489: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F(26),
  I1 => R1IN_2_2F(9),
  O => R1IN_2_ADD_1_AXB_9);
R1IN_2_ADD_1_AXB_10_Z5490: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F(27),
  I1 => R1IN_2_2F(10),
  O => R1IN_2_ADD_1_AXB_10);
R1IN_2_ADD_1_AXB_11_Z5491: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F(28),
  I1 => R1IN_2_2F(11),
  O => R1IN_2_ADD_1_AXB_11);
R1IN_2_ADD_1_AXB_12_Z5492: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F(29),
  I1 => R1IN_2_2F(12),
  O => R1IN_2_ADD_1_AXB_12);
R1IN_2_ADD_1_AXB_13_Z5493: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F(30),
  I1 => R1IN_2_2F(13),
  O => R1IN_2_ADD_1_AXB_13);
R1IN_2_ADD_1_AXB_14_Z5494: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F(31),
  I1 => R1IN_2_2F(14),
  O => R1IN_2_ADD_1_AXB_14);
R1IN_2_ADD_1_AXB_15_Z5495: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F(32),
  I1 => R1IN_2_2F(15),
  O => R1IN_2_ADD_1_AXB_15);
R1IN_2_ADD_1_AXB_16_Z5496: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2_1F(33),
  I1 => R1IN_2_2F(16),
  O => R1IN_2_ADD_1_AXB_16);
R1IN_2_ADD_1_AXB_17_Z5497: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(17),
  O => R1IN_2_ADD_1_AXB_17);
R1IN_2_ADD_1_AXB_18_Z5498: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(18),
  O => R1IN_2_ADD_1_AXB_18);
R1IN_2_ADD_1_AXB_19_Z5499: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(19),
  O => R1IN_2_ADD_1_AXB_19);
R1IN_2_ADD_1_AXB_20_Z5500: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(20),
  O => R1IN_2_ADD_1_AXB_20);
R1IN_2_ADD_1_AXB_21_Z5501: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(21),
  O => R1IN_2_ADD_1_AXB_21);
R1IN_2_ADD_1_AXB_22_Z5502: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(22),
  O => R1IN_2_ADD_1_AXB_22);
R1IN_2_ADD_1_AXB_23_Z5503: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(23),
  O => R1IN_2_ADD_1_AXB_23);
R1IN_2_ADD_1_AXB_24_Z5504: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(24),
  O => R1IN_2_ADD_1_AXB_24);
R1IN_2_ADD_1_AXB_25_Z5505: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(25),
  O => R1IN_2_ADD_1_AXB_25);
R1IN_2_ADD_1_AXB_26_Z5506: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(26),
  O => R1IN_2_ADD_1_AXB_26);
R1IN_2_ADD_1_AXB_27_Z5507: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(27),
  O => R1IN_2_ADD_1_AXB_27);
R1IN_2_ADD_1_AXB_28_Z5508: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(28),
  O => R1IN_2_ADD_1_AXB_28);
R1IN_2_ADD_1_AXB_29_Z5509: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(29),
  O => R1IN_2_ADD_1_AXB_29);
R1IN_2_ADD_1_AXB_30_Z5510: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(30),
  O => R1IN_2_ADD_1_AXB_30);
R1IN_2_ADD_1_AXB_31_Z5511: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(31),
  O => R1IN_2_ADD_1_AXB_31);
R1IN_2_ADD_1_AXB_32_Z5512: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(32),
  O => R1IN_2_ADD_1_AXB_32);
R1IN_2_ADD_1_AXB_33_Z5513: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(33),
  O => R1IN_2_ADD_1_AXB_33);
R1IN_2_ADD_1_AXB_34_Z5514: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(34),
  O => R1IN_2_ADD_1_AXB_34);
R1IN_2_ADD_1_AXB_35_Z5515: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(35),
  O => R1IN_2_ADD_1_AXB_35);
R1IN_2_ADD_1_AXB_36_Z5516: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(36),
  O => R1IN_2_ADD_1_AXB_36);
R1IN_2_ADD_1_AXB_37_Z5517: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(37),
  O => R1IN_2_ADD_1_AXB_37);
R1IN_2_ADD_1_AXB_38_Z5518: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(38),
  O => R1IN_2_ADD_1_AXB_38);
R1IN_2_ADD_1_AXB_39_Z5519: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(39),
  O => R1IN_2_ADD_1_AXB_39);
R1IN_2_ADD_1_AXB_40_Z5520: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(40),
  O => R1IN_2_ADD_1_AXB_40);
R1IN_2_ADD_1_AXB_41_Z5521: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(41),
  O => R1IN_2_ADD_1_AXB_41);
R1IN_2_ADD_1_AXB_42_Z5522: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(42),
  O => R1IN_2_ADD_1_AXB_42);
R1IN_4_4_ADD_2_AXB_1_Z5523: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F(18),
  I1 => R1IN_4_4_ADD_1F(1),
  O => R1IN_4_4_ADD_2_AXB_1);
R1IN_4_4_ADD_2_AXB_2_Z5524: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F(19),
  I1 => R1IN_4_4_ADD_1F(2),
  O => R1IN_4_4_ADD_2_AXB_2);
R1IN_4_4_ADD_2_AXB_3_Z5525: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F(20),
  I1 => R1IN_4_4_ADD_1F(3),
  O => R1IN_4_4_ADD_2_AXB_3);
R1IN_4_4_ADD_2_AXB_4_Z5526: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F(21),
  I1 => R1IN_4_4_ADD_1F(4),
  O => R1IN_4_4_ADD_2_AXB_4);
R1IN_4_4_ADD_2_AXB_5_Z5527: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F(22),
  I1 => R1IN_4_4_ADD_1F(5),
  O => R1IN_4_4_ADD_2_AXB_5);
R1IN_4_4_ADD_2_AXB_6_Z5528: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F(23),
  I1 => R1IN_4_4_ADD_1F(6),
  O => R1IN_4_4_ADD_2_AXB_6);
R1IN_4_4_ADD_2_AXB_7_Z5529: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F(24),
  I1 => R1IN_4_4_ADD_1F(7),
  O => R1IN_4_4_ADD_2_AXB_7);
R1IN_4_4_ADD_2_AXB_8_Z5530: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F(25),
  I1 => R1IN_4_4_ADD_1F(8),
  O => R1IN_4_4_ADD_2_AXB_8);
R1IN_4_4_ADD_2_AXB_9_Z5531: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F(26),
  I1 => R1IN_4_4_ADD_1F(9),
  O => R1IN_4_4_ADD_2_AXB_9);
R1IN_4_4_ADD_2_AXB_10_Z5532: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F(27),
  I1 => R1IN_4_4_ADD_1F(10),
  O => R1IN_4_4_ADD_2_AXB_10);
R1IN_4_4_ADD_2_AXB_11_Z5533: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F(28),
  I1 => R1IN_4_4_ADD_1F(11),
  O => R1IN_4_4_ADD_2_AXB_11);
R1IN_4_4_ADD_2_AXB_12_Z5534: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F(29),
  I1 => R1IN_4_4_ADD_1F(12),
  O => R1IN_4_4_ADD_2_AXB_12);
R1IN_4_4_ADD_2_AXB_13_Z5535: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F(30),
  I1 => R1IN_4_4_ADD_1F(13),
  O => R1IN_4_4_ADD_2_AXB_13);
R1IN_4_4_ADD_2_AXB_14_Z5536: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F(31),
  I1 => R1IN_4_4_ADD_1F(14),
  O => R1IN_4_4_ADD_2_AXB_14);
R1IN_4_4_ADD_2_AXB_15_Z5537: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F(32),
  I1 => R1IN_4_4_ADD_1F(15),
  O => R1IN_4_4_ADD_2_AXB_15);
R1IN_4_4_ADD_2_AXB_16_Z5538: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_1F(33),
  I1 => R1IN_4_4_ADD_1F(16),
  O => R1IN_4_4_ADD_2_AXB_16);
R1IN_4_4_ADD_2_AXB_17_Z5539: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_4F(0),
  I1 => R1IN_4_4_ADD_1F(17),
  O => R1IN_4_4_ADD_2_AXB_17);
R1IN_4_4_ADD_2_AXB_18_Z5540: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_4F(1),
  I1 => R1IN_4_4_ADD_1F(18),
  O => R1IN_4_4_ADD_2_AXB_18);
R1IN_4_4_ADD_2_AXB_19_Z5541: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_4F(2),
  I1 => R1IN_4_4_ADD_1F(19),
  O => R1IN_4_4_ADD_2_AXB_19);
R1IN_4_4_ADD_2_AXB_20_Z5542: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_4F(3),
  I1 => R1IN_4_4_ADD_1F(20),
  O => R1IN_4_4_ADD_2_AXB_20);
R1IN_4_4_ADD_2_AXB_21_Z5543: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_4F(4),
  I1 => R1IN_4_4_ADD_1F(21),
  O => R1IN_4_4_ADD_2_AXB_21);
R1IN_4_4_ADD_2_AXB_22_Z5544: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_4F(5),
  I1 => R1IN_4_4_ADD_1F(22),
  O => R1IN_4_4_ADD_2_AXB_22);
R1IN_4_4_ADD_2_AXB_23_Z5545: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_4F(6),
  I1 => R1IN_4_4_ADD_1F(23),
  O => R1IN_4_4_ADD_2_AXB_23);
R1IN_4_4_ADD_2_AXB_24_Z5546: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_4F(7),
  I1 => R1IN_4_4_ADD_1F(24),
  O => R1IN_4_4_ADD_2_AXB_24);
R1IN_4_4_ADD_2_AXB_25_Z5547: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_4F(8),
  I1 => R1IN_4_4_ADD_1F(25),
  O => R1IN_4_4_ADD_2_AXB_25);
R1IN_4_4_ADD_2_AXB_26_Z5548: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_4F(9),
  I1 => R1IN_4_4_ADD_1F(26),
  O => R1IN_4_4_ADD_2_AXB_26);
R1IN_4_4_ADD_2_AXB_27_Z5549: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_4F(10),
  I1 => R1IN_4_4_ADD_1F(27),
  O => R1IN_4_4_ADD_2_AXB_27);
R1IN_4_4_ADD_2_AXB_28_Z5550: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4_4F(11),
  O => R1IN_4_4_ADD_2_AXB_28);
R1IN_4_4_ADD_2_AXB_29_Z5551: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4_4F(12),
  O => R1IN_4_4_ADD_2_AXB_29);
R1IN_4_4_ADD_2_AXB_30_Z5552: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4_4F(13),
  O => R1IN_4_4_ADD_2_AXB_30);
R1IN_4_4_ADD_2_AXB_31_Z5553: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4_4F(14),
  O => R1IN_4_4_ADD_2_AXB_31);
R1IN_4_4_ADD_2_AXB_32_Z5554: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4_4F(15),
  O => R1IN_4_4_ADD_2_AXB_32);
R1IN_4_4_ADD_2_AXB_33_Z5555: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4_4F(16),
  O => R1IN_4_4_ADD_2_AXB_33);
R1IN_4_4_ADD_2_AXB_34_Z5556: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4_4F(17),
  O => R1IN_4_4_ADD_2_AXB_34);
R1IN_4_4_ADD_2_AXB_35_Z5557: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4_4F(18),
  O => R1IN_4_4_ADD_2_AXB_35);
R1IN_4_ADD_1_AXB_1_Z5558: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(1),
  I1 => R1IN_4_3F(1),
  O => R1IN_4_ADD_1_AXB_1);
R1IN_4_ADD_1_AXB_2_Z5559: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(2),
  I1 => R1IN_4_3F(2),
  O => R1IN_4_ADD_1_AXB_2);
R1IN_4_ADD_1_AXB_3_Z5560: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(3),
  I1 => R1IN_4_3F(3),
  O => R1IN_4_ADD_1_AXB_3);
R1IN_4_ADD_1_AXB_4_Z5561: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(4),
  I1 => R1IN_4_3F(4),
  O => R1IN_4_ADD_1_AXB_4);
R1IN_4_ADD_1_AXB_5_Z5562: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(5),
  I1 => R1IN_4_3F(5),
  O => R1IN_4_ADD_1_AXB_5);
R1IN_4_ADD_1_AXB_6_Z5563: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(6),
  I1 => R1IN_4_3F(6),
  O => R1IN_4_ADD_1_AXB_6);
R1IN_4_ADD_1_AXB_7_Z5564: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(7),
  I1 => R1IN_4_3F(7),
  O => R1IN_4_ADD_1_AXB_7);
R1IN_4_ADD_1_AXB_8_Z5565: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(8),
  I1 => R1IN_4_3F(8),
  O => R1IN_4_ADD_1_AXB_8);
R1IN_4_ADD_1_AXB_9_Z5566: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(9),
  I1 => R1IN_4_3F(9),
  O => R1IN_4_ADD_1_AXB_9);
R1IN_4_ADD_1_AXB_10_Z5567: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(10),
  I1 => R1IN_4_3F(10),
  O => R1IN_4_ADD_1_AXB_10);
R1IN_4_ADD_1_AXB_11_Z5568: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(11),
  I1 => R1IN_4_3F(11),
  O => R1IN_4_ADD_1_AXB_11);
R1IN_4_ADD_1_AXB_12_Z5569: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(12),
  I1 => R1IN_4_3F(12),
  O => R1IN_4_ADD_1_AXB_12);
R1IN_4_ADD_1_AXB_13_Z5570: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(13),
  I1 => R1IN_4_3F(13),
  O => R1IN_4_ADD_1_AXB_13);
R1IN_4_ADD_1_AXB_14_Z5571: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(14),
  I1 => R1IN_4_3F(14),
  O => R1IN_4_ADD_1_AXB_14);
R1IN_4_ADD_1_AXB_15_Z5572: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(15),
  I1 => R1IN_4_3F(15),
  O => R1IN_4_ADD_1_AXB_15);
R1IN_4_ADD_1_AXB_16_Z5573: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(16),
  I1 => R1IN_4_3F(16),
  O => R1IN_4_ADD_1_AXB_16);
R1IN_4_ADD_1_AXB_17_Z5574: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(17),
  I1 => R1IN_4_3F(17),
  O => R1IN_4_ADD_1_AXB_17);
R1IN_4_ADD_1_AXB_18_Z5575: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(18),
  I1 => R1IN_4_3F(18),
  O => R1IN_4_ADD_1_AXB_18);
R1IN_4_ADD_1_AXB_19_Z5576: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(19),
  I1 => R1IN_4_3F(19),
  O => R1IN_4_ADD_1_AXB_19);
R1IN_4_ADD_1_AXB_20_Z5577: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(20),
  I1 => R1IN_4_3F(20),
  O => R1IN_4_ADD_1_AXB_20);
R1IN_4_ADD_1_AXB_21_Z5578: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(21),
  I1 => R1IN_4_3F(21),
  O => R1IN_4_ADD_1_AXB_21);
R1IN_4_ADD_1_AXB_22_Z5579: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(22),
  I1 => R1IN_4_3F(22),
  O => R1IN_4_ADD_1_AXB_22);
R1IN_4_ADD_1_AXB_23_Z5580: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(23),
  I1 => R1IN_4_3F(23),
  O => R1IN_4_ADD_1_AXB_23);
R1IN_4_ADD_1_AXB_24_Z5581: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(24),
  I1 => R1IN_4_3F(24),
  O => R1IN_4_ADD_1_AXB_24);
R1IN_4_ADD_1_AXB_25_Z5582: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(25),
  I1 => R1IN_4_3F(25),
  O => R1IN_4_ADD_1_AXB_25);
R1IN_4_ADD_1_AXB_26_Z5583: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(26),
  I1 => R1IN_4_3F(26),
  O => R1IN_4_ADD_1_AXB_26);
R1IN_4_ADD_1_AXB_27_Z5584: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(27),
  I1 => R1IN_4_3F(27),
  O => R1IN_4_ADD_1_AXB_27);
R1IN_4_ADD_1_AXB_28_Z5585: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(28),
  I1 => R1IN_4_3F(28),
  O => R1IN_4_ADD_1_AXB_28);
R1IN_4_ADD_1_AXB_29_Z5586: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(29),
  I1 => R1IN_4_3F(29),
  O => R1IN_4_ADD_1_AXB_29);
R1IN_4_ADD_1_AXB_30_Z5587: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(30),
  I1 => R1IN_4_3F(30),
  O => R1IN_4_ADD_1_AXB_30);
R1IN_4_ADD_1_AXB_31_Z5588: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(31),
  I1 => R1IN_4_3F(31),
  O => R1IN_4_ADD_1_AXB_31);
R1IN_4_ADD_1_AXB_32_Z5589: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(32),
  I1 => R1IN_4_3F(32),
  O => R1IN_4_ADD_1_AXB_32);
R1IN_4_ADD_1_AXB_33_Z5590: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(33),
  I1 => R1IN_4_3F(33),
  O => R1IN_4_ADD_1_AXB_33);
R1IN_4_ADD_1_AXB_34_Z5591: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(34),
  I1 => R1IN_4_3F(34),
  O => R1IN_4_ADD_1_AXB_34);
R1IN_4_ADD_1_AXB_35_Z5592: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(35),
  I1 => R1IN_4_3F(35),
  O => R1IN_4_ADD_1_AXB_35);
R1IN_4_ADD_1_AXB_36_Z5593: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(36),
  I1 => R1IN_4_3F(36),
  O => R1IN_4_ADD_1_AXB_36);
R1IN_4_ADD_1_AXB_37_Z5594: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(37),
  I1 => R1IN_4_3F(37),
  O => R1IN_4_ADD_1_AXB_37);
R1IN_4_ADD_1_AXB_38_Z5595: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(38),
  I1 => R1IN_4_3F(38),
  O => R1IN_4_ADD_1_AXB_38);
R1IN_4_ADD_1_AXB_39_Z5596: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(39),
  I1 => R1IN_4_3F(39),
  O => R1IN_4_ADD_1_AXB_39);
R1IN_4_ADD_1_AXB_40_Z5597: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(40),
  I1 => R1IN_4_3F(40),
  O => R1IN_4_ADD_1_AXB_40);
R1IN_4_ADD_1_AXB_41_Z5598: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(41),
  I1 => R1IN_4_3F(41),
  O => R1IN_4_ADD_1_AXB_41);
R1IN_4_ADD_1_AXB_42_Z5599: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(42),
  I1 => R1IN_4_3F(42),
  O => R1IN_4_ADD_1_AXB_42);
R1IN_4_ADD_1_AXB_43_Z5600: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_2F(43),
  I1 => R1IN_4_3F(43),
  O => R1IN_4_ADD_1_AXB_43);
R1_PIPE_34: FDE port map (
    Q => NN_12,
    D => R1IN_4_2(0),
    C => CLK,
    CE => EN);
R1_PIPE_283: FDE port map (
    Q => R1IN_4_2F(1),
    D => R1IN_4_2(1),
    C => CLK,
    CE => EN);
R1_PIPE_284: FDE port map (
    Q => R1IN_4_2F(2),
    D => R1IN_4_2(2),
    C => CLK,
    CE => EN);
R1_PIPE_285: FDE port map (
    Q => R1IN_4_2F(3),
    D => R1IN_4_2(3),
    C => CLK,
    CE => EN);
R1_PIPE_286: FDE port map (
    Q => R1IN_4_2F(4),
    D => R1IN_4_2(4),
    C => CLK,
    CE => EN);
R1_PIPE_287: FDE port map (
    Q => R1IN_4_2F(5),
    D => R1IN_4_2(5),
    C => CLK,
    CE => EN);
R1_PIPE_288: FDE port map (
    Q => R1IN_4_2F(6),
    D => R1IN_4_2(6),
    C => CLK,
    CE => EN);
R1_PIPE_289: FDE port map (
    Q => R1IN_4_2F(7),
    D => R1IN_4_2(7),
    C => CLK,
    CE => EN);
R1_PIPE_290: FDE port map (
    Q => R1IN_4_2F(8),
    D => R1IN_4_2(8),
    C => CLK,
    CE => EN);
R1_PIPE_291: FDE port map (
    Q => R1IN_4_2F(9),
    D => R1IN_4_2(9),
    C => CLK,
    CE => EN);
R1_PIPE_292: FDE port map (
    Q => R1IN_4_2F(10),
    D => R1IN_4_2(10),
    C => CLK,
    CE => EN);
R1_PIPE_293: FDE port map (
    Q => R1IN_4_2F(11),
    D => R1IN_4_2(11),
    C => CLK,
    CE => EN);
R1_PIPE_294: FDE port map (
    Q => R1IN_4_2F(12),
    D => R1IN_4_2(12),
    C => CLK,
    CE => EN);
R1_PIPE_295: FDE port map (
    Q => R1IN_4_2F(13),
    D => R1IN_4_2(13),
    C => CLK,
    CE => EN);
R1_PIPE_296: FDE port map (
    Q => R1IN_4_2F(14),
    D => R1IN_4_2(14),
    C => CLK,
    CE => EN);
R1_PIPE_297: FDE port map (
    Q => R1IN_4_2F(15),
    D => R1IN_4_2(15),
    C => CLK,
    CE => EN);
R1_PIPE_298: FDE port map (
    Q => R1IN_4_2F(16),
    D => R1IN_4_2(16),
    C => CLK,
    CE => EN);
R1_PIPE_326: FDE port map (
    Q => R1IN_4_3F(0),
    D => R1IN_4_3(0),
    C => CLK,
    CE => EN);
R1_PIPE_327: FDE port map (
    Q => R1IN_4_3F(1),
    D => R1IN_4_3(1),
    C => CLK,
    CE => EN);
R1_PIPE_328: FDE port map (
    Q => R1IN_4_3F(2),
    D => R1IN_4_3(2),
    C => CLK,
    CE => EN);
R1_PIPE_329: FDE port map (
    Q => R1IN_4_3F(3),
    D => R1IN_4_3(3),
    C => CLK,
    CE => EN);
R1_PIPE_330: FDE port map (
    Q => R1IN_4_3F(4),
    D => R1IN_4_3(4),
    C => CLK,
    CE => EN);
R1_PIPE_331: FDE port map (
    Q => R1IN_4_3F(5),
    D => R1IN_4_3(5),
    C => CLK,
    CE => EN);
R1_PIPE_332: FDE port map (
    Q => R1IN_4_3F(6),
    D => R1IN_4_3(6),
    C => CLK,
    CE => EN);
R1_PIPE_333: FDE port map (
    Q => R1IN_4_3F(7),
    D => R1IN_4_3(7),
    C => CLK,
    CE => EN);
R1_PIPE_334: FDE port map (
    Q => R1IN_4_3F(8),
    D => R1IN_4_3(8),
    C => CLK,
    CE => EN);
R1_PIPE_335: FDE port map (
    Q => R1IN_4_3F(9),
    D => R1IN_4_3(9),
    C => CLK,
    CE => EN);
R1_PIPE_336: FDE port map (
    Q => R1IN_4_3F(10),
    D => R1IN_4_3(10),
    C => CLK,
    CE => EN);
R1_PIPE_337: FDE port map (
    Q => R1IN_4_3F(11),
    D => R1IN_4_3(11),
    C => CLK,
    CE => EN);
R1_PIPE_338: FDE port map (
    Q => R1IN_4_3F(12),
    D => R1IN_4_3(12),
    C => CLK,
    CE => EN);
R1_PIPE_339: FDE port map (
    Q => R1IN_4_3F(13),
    D => R1IN_4_3(13),
    C => CLK,
    CE => EN);
R1_PIPE_340: FDE port map (
    Q => R1IN_4_3F(14),
    D => R1IN_4_3(14),
    C => CLK,
    CE => EN);
R1_PIPE_341: FDE port map (
    Q => R1IN_4_3F(15),
    D => R1IN_4_3(15),
    C => CLK,
    CE => EN);
R1_PIPE_342: FDE port map (
    Q => R1IN_4_3F(16),
    D => R1IN_4_3(16),
    C => CLK,
    CE => EN);
R2_PIPE_17: FDE port map (
    Q => R1IN_4FF(0),
    D => R1IN_4F(0),
    C => CLK,
    CE => EN);
R2_PIPE_18: FDE port map (
    Q => R1IN_4FF(1),
    D => R1IN_4F(1),
    C => CLK,
    CE => EN);
R2_PIPE_19: FDE port map (
    Q => R1IN_4FF(2),
    D => R1IN_4F(2),
    C => CLK,
    CE => EN);
R2_PIPE_20: FDE port map (
    Q => R1IN_4FF(3),
    D => R1IN_4F(3),
    C => CLK,
    CE => EN);
R2_PIPE_21: FDE port map (
    Q => R1IN_4FF(4),
    D => R1IN_4F(4),
    C => CLK,
    CE => EN);
R2_PIPE_22: FDE port map (
    Q => R1IN_4FF(5),
    D => R1IN_4F(5),
    C => CLK,
    CE => EN);
R2_PIPE_23: FDE port map (
    Q => R1IN_4FF(6),
    D => R1IN_4F(6),
    C => CLK,
    CE => EN);
R2_PIPE_24: FDE port map (
    Q => R1IN_4FF(7),
    D => R1IN_4F(7),
    C => CLK,
    CE => EN);
R2_PIPE_25: FDE port map (
    Q => R1IN_4FF(8),
    D => R1IN_4F(8),
    C => CLK,
    CE => EN);
R2_PIPE_26: FDE port map (
    Q => R1IN_4FF(9),
    D => R1IN_4F(9),
    C => CLK,
    CE => EN);
R2_PIPE_27: FDE port map (
    Q => R1IN_4FF(10),
    D => R1IN_4F(10),
    C => CLK,
    CE => EN);
R2_PIPE_28: FDE port map (
    Q => R1IN_4FF(11),
    D => R1IN_4F(11),
    C => CLK,
    CE => EN);
R2_PIPE_29: FDE port map (
    Q => R1IN_4FF(12),
    D => R1IN_4F(12),
    C => CLK,
    CE => EN);
R2_PIPE_30: FDE port map (
    Q => R1IN_4FF(13),
    D => R1IN_4F(13),
    C => CLK,
    CE => EN);
R2_PIPE_31: FDE port map (
    Q => R1IN_4FF(14),
    D => R1IN_4F(14),
    C => CLK,
    CE => EN);
R2_PIPE_32: FDE port map (
    Q => R1IN_4FF(15),
    D => R1IN_4F(15),
    C => CLK,
    CE => EN);
R2_PIPE_33: FDE port map (
    Q => R1IN_4FF(16),
    D => R1IN_4F(16),
    C => CLK,
    CE => EN);
R2_PIPE_34: FDE port map (
    Q => R1IN_4F(17),
    D => R1IN_4(17),
    C => CLK,
    CE => EN);
R2_PIPE_35: FDE port map (
    Q => R1IN_4F(18),
    D => R1IN_4(18),
    C => CLK,
    CE => EN);
R2_PIPE_36: FDE port map (
    Q => R1IN_4F(19),
    D => R1IN_4(19),
    C => CLK,
    CE => EN);
R2_PIPE_37: FDE port map (
    Q => R1IN_4F(20),
    D => R1IN_4(20),
    C => CLK,
    CE => EN);
R2_PIPE_38: FDE port map (
    Q => R1IN_4F(21),
    D => R1IN_4(21),
    C => CLK,
    CE => EN);
R2_PIPE_39: FDE port map (
    Q => R1IN_4F(22),
    D => R1IN_4(22),
    C => CLK,
    CE => EN);
R2_PIPE_40: FDE port map (
    Q => R1IN_4F(23),
    D => R1IN_4(23),
    C => CLK,
    CE => EN);
R2_PIPE_41: FDE port map (
    Q => R1IN_4F(24),
    D => R1IN_4(24),
    C => CLK,
    CE => EN);
R2_PIPE_42: FDE port map (
    Q => R1IN_4F(25),
    D => R1IN_4(25),
    C => CLK,
    CE => EN);
R2_PIPE_43: FDE port map (
    Q => R1IN_4F(26),
    D => R1IN_4(26),
    C => CLK,
    CE => EN);
R2_PIPE_44: FDE port map (
    Q => R1IN_4F(27),
    D => R1IN_4(27),
    C => CLK,
    CE => EN);
R2_PIPE_45: FDE port map (
    Q => R1IN_4F(28),
    D => R1IN_4(28),
    C => CLK,
    CE => EN);
R2_PIPE_46: FDE port map (
    Q => R1IN_4F(29),
    D => R1IN_4(29),
    C => CLK,
    CE => EN);
R2_PIPE_47: FDE port map (
    Q => R1IN_4F(30),
    D => R1IN_4(30),
    C => CLK,
    CE => EN);
R2_PIPE_48: FDE port map (
    Q => R1IN_4F(31),
    D => R1IN_4(31),
    C => CLK,
    CE => EN);
R2_PIPE_49: FDE port map (
    Q => R1IN_4F(32),
    D => R1IN_4(32),
    C => CLK,
    CE => EN);
R2_PIPE_50: FDE port map (
    Q => R1IN_4F(33),
    D => R1IN_4(33),
    C => CLK,
    CE => EN);
R2_PIPE_51: FDE port map (
    Q => R1IN_4F(34),
    D => R1IN_4(34),
    C => CLK,
    CE => EN);
R2_PIPE_52: FDE port map (
    Q => R1IN_4F(35),
    D => R1IN_4(35),
    C => CLK,
    CE => EN);
R2_PIPE_53: FDE port map (
    Q => R1IN_4F(36),
    D => R1IN_4(36),
    C => CLK,
    CE => EN);
R2_PIPE_54: FDE port map (
    Q => R1IN_4F(37),
    D => R1IN_4(37),
    C => CLK,
    CE => EN);
R2_PIPE_55: FDE port map (
    Q => R1IN_4F(38),
    D => R1IN_4(38),
    C => CLK,
    CE => EN);
R2_PIPE_56: FDE port map (
    Q => R1IN_4F(39),
    D => R1IN_4(39),
    C => CLK,
    CE => EN);
R2_PIPE_57: FDE port map (
    Q => R1IN_4F(40),
    D => R1IN_4(40),
    C => CLK,
    CE => EN);
R2_PIPE_58: FDE port map (
    Q => R1IN_4F(41),
    D => R1IN_4(41),
    C => CLK,
    CE => EN);
R2_PIPE_59: FDE port map (
    Q => R1IN_4F(42),
    D => R1IN_4(42),
    C => CLK,
    CE => EN);
R2_PIPE_60: FDE port map (
    Q => R1IN_4F(43),
    D => R1IN_4(43),
    C => CLK,
    CE => EN);
R2_PIPE_61: FDE port map (
    Q => R1IN_4F(44),
    D => R1IN_4(44),
    C => CLK,
    CE => EN);
R2_PIPE_62: FDE port map (
    Q => R1IN_4F(45),
    D => R1IN_4(45),
    C => CLK,
    CE => EN);
R2_PIPE_63: FDE port map (
    Q => R1IN_4F(46),
    D => R1IN_4(46),
    C => CLK,
    CE => EN);
R2_PIPE_64: FDE port map (
    Q => R1IN_4F(47),
    D => R1IN_4(47),
    C => CLK,
    CE => EN);
R2_PIPE_65: FDE port map (
    Q => R1IN_4F(48),
    D => R1IN_4(48),
    C => CLK,
    CE => EN);
R2_PIPE_66: FDE port map (
    Q => R1IN_4F(49),
    D => R1IN_4(49),
    C => CLK,
    CE => EN);
R2_PIPE_67: FDE port map (
    Q => R1IN_4F(50),
    D => R1IN_4(50),
    C => CLK,
    CE => EN);
R2_PIPE_68: FDE port map (
    Q => R1IN_4F(51),
    D => R1IN_4(51),
    C => CLK,
    CE => EN);
R2_PIPE_69: FDE port map (
    Q => R1IN_4F(52),
    D => R1IN_4(52),
    C => CLK,
    CE => EN);
R2_PIPE_105: FDE port map (
    Q => R1IN_ADD_1FF(0),
    D => R1IN_ADD_1(0),
    C => CLK,
    CE => EN);
R2_PIPE_106: FDE port map (
    Q => R1IN_ADD_1FF(1),
    D => R1IN_ADD_1(1),
    C => CLK,
    CE => EN);
R2_PIPE_107: FDE port map (
    Q => R1IN_ADD_1FF(2),
    D => R1IN_ADD_1(2),
    C => CLK,
    CE => EN);
R2_PIPE_108: FDE port map (
    Q => R1IN_ADD_1FF(3),
    D => R1IN_ADD_1(3),
    C => CLK,
    CE => EN);
R2_PIPE_109: FDE port map (
    Q => R1IN_ADD_1FF(4),
    D => R1IN_ADD_1(4),
    C => CLK,
    CE => EN);
R2_PIPE_110: FDE port map (
    Q => R1IN_ADD_1FF(5),
    D => R1IN_ADD_1(5),
    C => CLK,
    CE => EN);
R2_PIPE_111: FDE port map (
    Q => R1IN_ADD_1FF(6),
    D => R1IN_ADD_1(6),
    C => CLK,
    CE => EN);
R2_PIPE_112: FDE port map (
    Q => R1IN_ADD_1FF(7),
    D => R1IN_ADD_1(7),
    C => CLK,
    CE => EN);
R2_PIPE_113: FDE port map (
    Q => R1IN_ADD_1FF(8),
    D => R1IN_ADD_1(8),
    C => CLK,
    CE => EN);
R2_PIPE_114: FDE port map (
    Q => R1IN_ADD_1FF(9),
    D => R1IN_ADD_1(9),
    C => CLK,
    CE => EN);
R2_PIPE_115: FDE port map (
    Q => R1IN_ADD_1FF(10),
    D => R1IN_ADD_1(10),
    C => CLK,
    CE => EN);
R2_PIPE_116: FDE port map (
    Q => R1IN_ADD_1FF(11),
    D => R1IN_ADD_1(11),
    C => CLK,
    CE => EN);
R2_PIPE_117: FDE port map (
    Q => R1IN_ADD_1FF(12),
    D => R1IN_ADD_1(12),
    C => CLK,
    CE => EN);
R2_PIPE_118: FDE port map (
    Q => R1IN_ADD_1FF(13),
    D => R1IN_ADD_1(13),
    C => CLK,
    CE => EN);
R2_PIPE_119: FDE port map (
    Q => R1IN_ADD_1FF(14),
    D => R1IN_ADD_1(14),
    C => CLK,
    CE => EN);
R2_PIPE_120: FDE port map (
    Q => R1IN_ADD_1FF(15),
    D => R1IN_ADD_1(15),
    C => CLK,
    CE => EN);
R2_PIPE_121: FDE port map (
    Q => R1IN_ADD_1FF(16),
    D => R1IN_ADD_1(16),
    C => CLK,
    CE => EN);
R2_PIPE_122: FDE port map (
    Q => R1IN_ADD_1FF(17),
    D => R1IN_ADD_1(17),
    C => CLK,
    CE => EN);
R2_PIPE_123: FDE port map (
    Q => R1IN_ADD_1FF(18),
    D => R1IN_ADD_1(18),
    C => CLK,
    CE => EN);
R2_PIPE_124: FDE port map (
    Q => R1IN_ADD_1FF(19),
    D => R1IN_ADD_1(19),
    C => CLK,
    CE => EN);
R2_PIPE_125: FDE port map (
    Q => R1IN_ADD_1FF(20),
    D => R1IN_ADD_1(20),
    C => CLK,
    CE => EN);
R2_PIPE_126: FDE port map (
    Q => R1IN_ADD_1FF(21),
    D => R1IN_ADD_1(21),
    C => CLK,
    CE => EN);
R2_PIPE_127: FDE port map (
    Q => R1IN_ADD_1FF(22),
    D => R1IN_ADD_1(22),
    C => CLK,
    CE => EN);
R2_PIPE_128: FDE port map (
    Q => R1IN_ADD_1FF(23),
    D => R1IN_ADD_1(23),
    C => CLK,
    CE => EN);
R2_PIPE_129: FDE port map (
    Q => R1IN_ADD_1FF(24),
    D => R1IN_ADD_1(24),
    C => CLK,
    CE => EN);
R2_PIPE_130: FDE port map (
    Q => R1IN_ADD_1FF(25),
    D => R1IN_ADD_1(25),
    C => CLK,
    CE => EN);
R2_PIPE_131: FDE port map (
    Q => R1IN_ADD_1FF(26),
    D => R1IN_ADD_1(26),
    C => CLK,
    CE => EN);
R2_PIPE_132: FDE port map (
    Q => R1IN_ADD_1FF(27),
    D => R1IN_ADD_1(27),
    C => CLK,
    CE => EN);
R2_PIPE_133: FDE port map (
    Q => R1IN_ADD_1FF(28),
    D => R1IN_ADD_1(28),
    C => CLK,
    CE => EN);
R2_PIPE_134: FDE port map (
    Q => R1IN_ADD_1FF(29),
    D => R1IN_ADD_1(29),
    C => CLK,
    CE => EN);
R2_PIPE_135: FDE port map (
    Q => R1IN_ADD_1FF(30),
    D => R1IN_ADD_1(30),
    C => CLK,
    CE => EN);
R2_PIPE_136: FDE port map (
    Q => R1IN_ADD_1FF(31),
    D => R1IN_ADD_1(31),
    C => CLK,
    CE => EN);
R2_PIPE_137: FDE port map (
    Q => R1IN_ADD_1FF(32),
    D => R1IN_ADD_1(32),
    C => CLK,
    CE => EN);
R1_PIPE_105: FDE port map (
    Q => R1IN_2_ADD_1,
    D => R1IN_2_2(0),
    C => CLK,
    CE => EN);
R1_PIPE_589: FDE port map (
    Q => R1IN_2_2F(1),
    D => R1IN_2_2(1),
    C => CLK,
    CE => EN);
R1_PIPE_590: FDE port map (
    Q => R1IN_2_2F(2),
    D => R1IN_2_2(2),
    C => CLK,
    CE => EN);
R1_PIPE_591: FDE port map (
    Q => R1IN_2_2F(3),
    D => R1IN_2_2(3),
    C => CLK,
    CE => EN);
R1_PIPE_592: FDE port map (
    Q => R1IN_2_2F(4),
    D => R1IN_2_2(4),
    C => CLK,
    CE => EN);
R1_PIPE_593: FDE port map (
    Q => R1IN_2_2F(5),
    D => R1IN_2_2(5),
    C => CLK,
    CE => EN);
R1_PIPE_594: FDE port map (
    Q => R1IN_2_2F(6),
    D => R1IN_2_2(6),
    C => CLK,
    CE => EN);
R1_PIPE_595: FDE port map (
    Q => R1IN_2_2F(7),
    D => R1IN_2_2(7),
    C => CLK,
    CE => EN);
R1_PIPE_596: FDE port map (
    Q => R1IN_2_2F(8),
    D => R1IN_2_2(8),
    C => CLK,
    CE => EN);
R1_PIPE_597: FDE port map (
    Q => R1IN_2_2F(9),
    D => R1IN_2_2(9),
    C => CLK,
    CE => EN);
R1_PIPE_598: FDE port map (
    Q => R1IN_2_2F(10),
    D => R1IN_2_2(10),
    C => CLK,
    CE => EN);
R1_PIPE_599: FDE port map (
    Q => R1IN_2_2F(11),
    D => R1IN_2_2(11),
    C => CLK,
    CE => EN);
R1_PIPE_600: FDE port map (
    Q => R1IN_2_2F(12),
    D => R1IN_2_2(12),
    C => CLK,
    CE => EN);
R1_PIPE_601: FDE port map (
    Q => R1IN_2_2F(13),
    D => R1IN_2_2(13),
    C => CLK,
    CE => EN);
R1_PIPE_602: FDE port map (
    Q => R1IN_2_2F(14),
    D => R1IN_2_2(14),
    C => CLK,
    CE => EN);
R1_PIPE_603: FDE port map (
    Q => R1IN_2_2F(15),
    D => R1IN_2_2(15),
    C => CLK,
    CE => EN);
R1_PIPE_604: FDE port map (
    Q => R1IN_2_2F(16),
    D => R1IN_2_2(16),
    C => CLK,
    CE => EN);
R1_PIPE_484: FDE port map (
    Q => R1IN_3_ADD_1,
    D => R1IN_3_2(0),
    C => CLK,
    CE => EN);
R1_PIPE_649: FDE port map (
    Q => R1IN_3_2F(1),
    D => R1IN_3_2(1),
    C => CLK,
    CE => EN);
R1_PIPE_650: FDE port map (
    Q => R1IN_3_2F(2),
    D => R1IN_3_2(2),
    C => CLK,
    CE => EN);
R1_PIPE_651: FDE port map (
    Q => R1IN_3_2F(3),
    D => R1IN_3_2(3),
    C => CLK,
    CE => EN);
R1_PIPE_652: FDE port map (
    Q => R1IN_3_2F(4),
    D => R1IN_3_2(4),
    C => CLK,
    CE => EN);
R1_PIPE_653: FDE port map (
    Q => R1IN_3_2F(5),
    D => R1IN_3_2(5),
    C => CLK,
    CE => EN);
R1_PIPE_654: FDE port map (
    Q => R1IN_3_2F(6),
    D => R1IN_3_2(6),
    C => CLK,
    CE => EN);
R1_PIPE_655: FDE port map (
    Q => R1IN_3_2F(7),
    D => R1IN_3_2(7),
    C => CLK,
    CE => EN);
R1_PIPE_656: FDE port map (
    Q => R1IN_3_2F(8),
    D => R1IN_3_2(8),
    C => CLK,
    CE => EN);
R1_PIPE_657: FDE port map (
    Q => R1IN_3_2F(9),
    D => R1IN_3_2(9),
    C => CLK,
    CE => EN);
R1_PIPE_658: FDE port map (
    Q => R1IN_3_2F(10),
    D => R1IN_3_2(10),
    C => CLK,
    CE => EN);
R1_PIPE_659: FDE port map (
    Q => R1IN_3_2F(11),
    D => R1IN_3_2(11),
    C => CLK,
    CE => EN);
R1_PIPE_660: FDE port map (
    Q => R1IN_3_2F(12),
    D => R1IN_3_2(12),
    C => CLK,
    CE => EN);
R1_PIPE_661: FDE port map (
    Q => R1IN_3_2F(13),
    D => R1IN_3_2(13),
    C => CLK,
    CE => EN);
R1_PIPE_662: FDE port map (
    Q => R1IN_3_2F(14),
    D => R1IN_3_2(14),
    C => CLK,
    CE => EN);
R1_PIPE_663: FDE port map (
    Q => R1IN_3_2F(15),
    D => R1IN_3_2(15),
    C => CLK,
    CE => EN);
R1_PIPE_664: FDE port map (
    Q => R1IN_3_2F(16),
    D => R1IN_3_2(16),
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_103_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_0,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_102_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_1,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_101_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_2,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_100_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_3,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_99_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_4,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_98_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_5,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_97_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_6,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_96_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_7,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_95_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_8,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_94_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_9,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_93_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_10,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_92_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_11,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_91_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_12,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_90_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_13,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_89_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_14,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_88_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_15,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_87_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_16,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_86_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_17,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_85_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_18,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_84_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_19,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_83_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_20,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_82_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_21,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_81_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_22,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_80_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_23,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_79_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_24,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_78_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_25,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_77_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_26,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_76_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_27,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_75_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_28,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_74_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_29,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_157_RET_Z5786: FDE port map (
    Q => R2_PIPE_157_RET,
    D => N_1577,
    C => CLK,
    CE => EN);
R2_PIPE_157_RET_1_Z5787: FDE port map (
    Q => R2_PIPE_157_RET_1,
    D => N_1913,
    C => CLK,
    CE => EN);
R2_PIPE_157_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_73_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_30,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_156_RET_Z5790: FDE port map (
    Q => R2_PIPE_156_RET,
    D => N_1575,
    C => CLK,
    CE => EN);
R2_PIPE_156_RET_1_Z5791: FDE port map (
    Q => R2_PIPE_156_RET_1,
    D => N_1912,
    C => CLK,
    CE => EN);
R2_PIPE_156_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_0,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_72_RET_2: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_31,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
R2_PIPE_155_RET_Z5794: FDE port map (
    Q => R2_PIPE_155_RET,
    D => N_1573,
    C => CLK,
    CE => EN);
R2_PIPE_155_RET_1_Z5795: FDE port map (
    Q => R2_PIPE_155_RET_1,
    D => N_1911,
    C => CLK,
    CE => EN);
R2_PIPE_155_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_1,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_154_RET_Z5797: FDE port map (
    Q => R2_PIPE_154_RET,
    D => N_1571,
    C => CLK,
    CE => EN);
R2_PIPE_154_RET_1_Z5798: FDE port map (
    Q => R2_PIPE_154_RET_1,
    D => N_1910,
    C => CLK,
    CE => EN);
R2_PIPE_154_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_2,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_153_RET_Z5800: FDE port map (
    Q => R2_PIPE_153_RET,
    D => N_1569,
    C => CLK,
    CE => EN);
R2_PIPE_153_RET_1_Z5801: FDE port map (
    Q => R2_PIPE_153_RET_1,
    D => N_1909,
    C => CLK,
    CE => EN);
R2_PIPE_153_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_3,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_152_RET_Z5803: FDE port map (
    Q => R2_PIPE_152_RET,
    D => N_1567,
    C => CLK,
    CE => EN);
R2_PIPE_152_RET_1_Z5804: FDE port map (
    Q => R2_PIPE_152_RET_1,
    D => N_1908,
    C => CLK,
    CE => EN);
R2_PIPE_152_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_4,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_151_RET_Z5806: FDE port map (
    Q => R2_PIPE_151_RET,
    D => N_1565,
    C => CLK,
    CE => EN);
R2_PIPE_151_RET_1_Z5807: FDE port map (
    Q => R2_PIPE_151_RET_1,
    D => N_1907,
    C => CLK,
    CE => EN);
R2_PIPE_151_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_5,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_150_RET_Z5809: FDE port map (
    Q => R2_PIPE_150_RET,
    D => N_1563,
    C => CLK,
    CE => EN);
R2_PIPE_150_RET_1_Z5810: FDE port map (
    Q => R2_PIPE_150_RET_1,
    D => N_1906,
    C => CLK,
    CE => EN);
R2_PIPE_150_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_6,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_149_RET_Z5812: FDE port map (
    Q => R2_PIPE_149_RET,
    D => N_1561,
    C => CLK,
    CE => EN);
R2_PIPE_149_RET_1_Z5813: FDE port map (
    Q => R2_PIPE_149_RET_1,
    D => N_1905,
    C => CLK,
    CE => EN);
R2_PIPE_149_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_7,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_148_RET_Z5815: FDE port map (
    Q => R2_PIPE_148_RET,
    D => N_1559,
    C => CLK,
    CE => EN);
R2_PIPE_148_RET_1_Z5816: FDE port map (
    Q => R2_PIPE_148_RET_1,
    D => N_1904,
    C => CLK,
    CE => EN);
R2_PIPE_148_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_8,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_147_RET_Z5818: FDE port map (
    Q => R2_PIPE_147_RET,
    D => N_1557,
    C => CLK,
    CE => EN);
R2_PIPE_147_RET_1_Z5819: FDE port map (
    Q => R2_PIPE_147_RET_1,
    D => N_1903,
    C => CLK,
    CE => EN);
R2_PIPE_147_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_9,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_146_RET_Z5821: FDE port map (
    Q => R2_PIPE_146_RET,
    D => N_1555,
    C => CLK,
    CE => EN);
R2_PIPE_146_RET_1_Z5822: FDE port map (
    Q => R2_PIPE_146_RET_1,
    D => N_1902,
    C => CLK,
    CE => EN);
R2_PIPE_146_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_10,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_145_RET_Z5824: FDE port map (
    Q => R2_PIPE_145_RET,
    D => N_1553,
    C => CLK,
    CE => EN);
R2_PIPE_145_RET_1_Z5825: FDE port map (
    Q => R2_PIPE_145_RET_1,
    D => N_1901,
    C => CLK,
    CE => EN);
R2_PIPE_145_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_11,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_144_RET_Z5827: FDE port map (
    Q => R2_PIPE_144_RET,
    D => N_1551,
    C => CLK,
    CE => EN);
R2_PIPE_144_RET_1_Z5828: FDE port map (
    Q => R2_PIPE_144_RET_1,
    D => N_1900,
    C => CLK,
    CE => EN);
R2_PIPE_144_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_12,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_143_RET_Z5830: FDE port map (
    Q => R2_PIPE_143_RET,
    D => N_1549,
    C => CLK,
    CE => EN);
R2_PIPE_143_RET_1_Z5831: FDE port map (
    Q => R2_PIPE_143_RET_1,
    D => N_1899,
    C => CLK,
    CE => EN);
R2_PIPE_143_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_13,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_142_RET_Z5833: FDE port map (
    Q => R2_PIPE_142_RET,
    D => N_1547,
    C => CLK,
    CE => EN);
R2_PIPE_142_RET_1_Z5834: FDE port map (
    Q => R2_PIPE_142_RET_1,
    D => N_1898,
    C => CLK,
    CE => EN);
R2_PIPE_142_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_14,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_141_RET_Z5836: FDE port map (
    Q => R2_PIPE_141_RET,
    D => N_1545,
    C => CLK,
    CE => EN);
R2_PIPE_141_RET_1_Z5837: FDE port map (
    Q => R2_PIPE_141_RET_1,
    D => N_1897,
    C => CLK,
    CE => EN);
R2_PIPE_141_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_15,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_140_RET_Z5839: FDE port map (
    Q => R2_PIPE_140_RET,
    D => N_1543,
    C => CLK,
    CE => EN);
R2_PIPE_140_RET_1_Z5840: FDE port map (
    Q => R2_PIPE_140_RET_1,
    D => N_1896,
    C => CLK,
    CE => EN);
R2_PIPE_140_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_16,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_139_RET_Z5842: FDE port map (
    Q => R2_PIPE_139_RET,
    D => N_1541,
    C => CLK,
    CE => EN);
R2_PIPE_139_RET_1_Z5843: FDE port map (
    Q => R2_PIPE_139_RET_1,
    D => N_1895,
    C => CLK,
    CE => EN);
R2_PIPE_139_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_17,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_138_RET_Z5845: FDE port map (
    Q => R2_PIPE_138_RET,
    D => N_1539,
    C => CLK,
    CE => EN);
R2_PIPE_138_RET_1_Z5846: FDE port map (
    Q => R2_PIPE_138_RET_1,
    D => N_1894,
    C => CLK,
    CE => EN);
R2_PIPE_138_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_18,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_3: FDE port map (
    Q => R1IN_4_ADD_2_0_CRY_35_RETO_32,
    D => R1IN_4_ADD_2_0_CRY_35,
    C => CLK,
    CE => EN);
\R1IN_3_1[0]\: FDE port map (
    Q => R1IN_3F(0),
    D => R1IN_3F_0(0),
    C => CLK,
    CE => EN);
\R1IN_3_1[1]\: FDE port map (
    Q => R1IN_3F(1),
    D => R1IN_3F_0(1),
    C => CLK,
    CE => EN);
\R1IN_3_1[2]\: FDE port map (
    Q => R1IN_3F(2),
    D => R1IN_3F_0(2),
    C => CLK,
    CE => EN);
\R1IN_3_1[3]\: FDE port map (
    Q => R1IN_3F(3),
    D => R1IN_3F_0(3),
    C => CLK,
    CE => EN);
\R1IN_3_1[4]\: FDE port map (
    Q => R1IN_3F(4),
    D => R1IN_3F_0(4),
    C => CLK,
    CE => EN);
\R1IN_3_1[5]\: FDE port map (
    Q => R1IN_3F(5),
    D => R1IN_3F_0(5),
    C => CLK,
    CE => EN);
\R1IN_3_1[6]\: FDE port map (
    Q => R1IN_3F(6),
    D => R1IN_3F_0(6),
    C => CLK,
    CE => EN);
\R1IN_3_1[7]\: FDE port map (
    Q => R1IN_3F(7),
    D => R1IN_3F_0(7),
    C => CLK,
    CE => EN);
\R1IN_3_1[8]\: FDE port map (
    Q => R1IN_3F(8),
    D => R1IN_3F_0(8),
    C => CLK,
    CE => EN);
\R1IN_3_1[9]\: FDE port map (
    Q => R1IN_3F(9),
    D => R1IN_3F_0(9),
    C => CLK,
    CE => EN);
\R1IN_3_1[10]\: FDE port map (
    Q => R1IN_3F(10),
    D => R1IN_3F_0(10),
    C => CLK,
    CE => EN);
\R1IN_3_1[11]\: FDE port map (
    Q => R1IN_3F(11),
    D => R1IN_3F_0(11),
    C => CLK,
    CE => EN);
\R1IN_3_1[12]\: FDE port map (
    Q => R1IN_3F(12),
    D => R1IN_3F_0(12),
    C => CLK,
    CE => EN);
\R1IN_3_1[13]\: FDE port map (
    Q => R1IN_3F(13),
    D => R1IN_3F_0(13),
    C => CLK,
    CE => EN);
\R1IN_3_1[14]\: FDE port map (
    Q => R1IN_3F(14),
    D => R1IN_3F_0(14),
    C => CLK,
    CE => EN);
\R1IN_3_1[15]\: FDE port map (
    Q => R1IN_3F(15),
    D => R1IN_3F_0(15),
    C => CLK,
    CE => EN);
\R1IN_3_1[16]\: FDE port map (
    Q => R1IN_3F(16),
    D => R1IN_3F_0(16),
    C => CLK,
    CE => EN);
\R1IN_3_1[17]\: FDE port map (
    Q => R1IN_3_1F(17),
    D => R1IN_3_1F_0(17),
    C => CLK,
    CE => EN);
\R1IN_3_1[18]\: FDE port map (
    Q => R1IN_3_1F(18),
    D => R1IN_3_1F_0(18),
    C => CLK,
    CE => EN);
\R1IN_3_1[19]\: FDE port map (
    Q => R1IN_3_1F(19),
    D => R1IN_3_1F_0(19),
    C => CLK,
    CE => EN);
\R1IN_3_1[20]\: FDE port map (
    Q => R1IN_3_1F(20),
    D => R1IN_3_1F_0(20),
    C => CLK,
    CE => EN);
\R1IN_3_1[21]\: FDE port map (
    Q => R1IN_3_1F(21),
    D => R1IN_3_1F_0(21),
    C => CLK,
    CE => EN);
\R1IN_3_1[22]\: FDE port map (
    Q => R1IN_3_1F(22),
    D => R1IN_3_1F_0(22),
    C => CLK,
    CE => EN);
\R1IN_3_1[23]\: FDE port map (
    Q => R1IN_3_1F(23),
    D => R1IN_3_1F_0(23),
    C => CLK,
    CE => EN);
\R1IN_3_1[24]\: FDE port map (
    Q => R1IN_3_1F(24),
    D => R1IN_3_1F_0(24),
    C => CLK,
    CE => EN);
\R1IN_3_1[25]\: FDE port map (
    Q => R1IN_3_1F(25),
    D => R1IN_3_1F_0(25),
    C => CLK,
    CE => EN);
\R1IN_3_1[26]\: FDE port map (
    Q => R1IN_3_1F(26),
    D => R1IN_3_1F_0(26),
    C => CLK,
    CE => EN);
\R1IN_3_1[27]\: FDE port map (
    Q => R1IN_3_1F(27),
    D => R1IN_3_1F_0(27),
    C => CLK,
    CE => EN);
\R1IN_3_1[28]\: FDE port map (
    Q => R1IN_3_1F(28),
    D => R1IN_3_1F_0(28),
    C => CLK,
    CE => EN);
\R1IN_3_1[29]\: FDE port map (
    Q => R1IN_3_1F(29),
    D => R1IN_3_1F_0(29),
    C => CLK,
    CE => EN);
\R1IN_3_1[30]\: FDE port map (
    Q => R1IN_3_1F(30),
    D => R1IN_3_1F_0(30),
    C => CLK,
    CE => EN);
\R1IN_3_1[31]\: FDE port map (
    Q => R1IN_3_1F(31),
    D => R1IN_3_1F_0(31),
    C => CLK,
    CE => EN);
\R1IN_3_1[32]\: FDE port map (
    Q => R1IN_3_1F(32),
    D => R1IN_3_1F_0(32),
    C => CLK,
    CE => EN);
\R1IN_3_1[33]\: FDE port map (
    Q => R1IN_3_1F(33),
    D => R1IN_3_1F_0(33),
    C => CLK,
    CE => EN);
\R1IN_2_1[0]\: FDE port map (
    Q => R1IN_2F(0),
    D => R1IN_2F_0(0),
    C => CLK,
    CE => EN);
\R1IN_2_1[1]\: FDE port map (
    Q => R1IN_2F(1),
    D => R1IN_2F_0(1),
    C => CLK,
    CE => EN);
\R1IN_2_1[2]\: FDE port map (
    Q => R1IN_2F(2),
    D => R1IN_2F_0(2),
    C => CLK,
    CE => EN);
\R1IN_2_1[3]\: FDE port map (
    Q => R1IN_2F(3),
    D => R1IN_2F_0(3),
    C => CLK,
    CE => EN);
\R1IN_2_1[4]\: FDE port map (
    Q => R1IN_2F(4),
    D => R1IN_2F_0(4),
    C => CLK,
    CE => EN);
\R1IN_2_1[5]\: FDE port map (
    Q => R1IN_2F(5),
    D => R1IN_2F_0(5),
    C => CLK,
    CE => EN);
\R1IN_2_1[6]\: FDE port map (
    Q => R1IN_2F(6),
    D => R1IN_2F_0(6),
    C => CLK,
    CE => EN);
\R1IN_2_1[7]\: FDE port map (
    Q => R1IN_2F(7),
    D => R1IN_2F_0(7),
    C => CLK,
    CE => EN);
\R1IN_2_1[8]\: FDE port map (
    Q => R1IN_2F(8),
    D => R1IN_2F_0(8),
    C => CLK,
    CE => EN);
\R1IN_2_1[9]\: FDE port map (
    Q => R1IN_2F(9),
    D => R1IN_2F_0(9),
    C => CLK,
    CE => EN);
\R1IN_2_1[10]\: FDE port map (
    Q => R1IN_2F(10),
    D => R1IN_2F_0(10),
    C => CLK,
    CE => EN);
\R1IN_2_1[11]\: FDE port map (
    Q => R1IN_2F(11),
    D => R1IN_2F_0(11),
    C => CLK,
    CE => EN);
\R1IN_2_1[12]\: FDE port map (
    Q => R1IN_2F(12),
    D => R1IN_2F_0(12),
    C => CLK,
    CE => EN);
\R1IN_2_1[13]\: FDE port map (
    Q => R1IN_2F(13),
    D => R1IN_2F_0(13),
    C => CLK,
    CE => EN);
\R1IN_2_1[14]\: FDE port map (
    Q => R1IN_2F(14),
    D => R1IN_2F_0(14),
    C => CLK,
    CE => EN);
\R1IN_2_1[15]\: FDE port map (
    Q => R1IN_2F(15),
    D => R1IN_2F_0(15),
    C => CLK,
    CE => EN);
\R1IN_2_1[16]\: FDE port map (
    Q => R1IN_2F(16),
    D => R1IN_2F_0(16),
    C => CLK,
    CE => EN);
\R1IN_2_1[17]\: FDE port map (
    Q => R1IN_2_1F(17),
    D => R1IN_2_1F_0(17),
    C => CLK,
    CE => EN);
\R1IN_2_1[18]\: FDE port map (
    Q => R1IN_2_1F(18),
    D => R1IN_2_1F_0(18),
    C => CLK,
    CE => EN);
\R1IN_2_1[19]\: FDE port map (
    Q => R1IN_2_1F(19),
    D => R1IN_2_1F_0(19),
    C => CLK,
    CE => EN);
\R1IN_2_1[20]\: FDE port map (
    Q => R1IN_2_1F(20),
    D => R1IN_2_1F_0(20),
    C => CLK,
    CE => EN);
\R1IN_2_1[21]\: FDE port map (
    Q => R1IN_2_1F(21),
    D => R1IN_2_1F_0(21),
    C => CLK,
    CE => EN);
\R1IN_2_1[22]\: FDE port map (
    Q => R1IN_2_1F(22),
    D => R1IN_2_1F_0(22),
    C => CLK,
    CE => EN);
\R1IN_2_1[23]\: FDE port map (
    Q => R1IN_2_1F(23),
    D => R1IN_2_1F_0(23),
    C => CLK,
    CE => EN);
\R1IN_2_1[24]\: FDE port map (
    Q => R1IN_2_1F(24),
    D => R1IN_2_1F_0(24),
    C => CLK,
    CE => EN);
\R1IN_2_1[25]\: FDE port map (
    Q => R1IN_2_1F(25),
    D => R1IN_2_1F_0(25),
    C => CLK,
    CE => EN);
\R1IN_2_1[26]\: FDE port map (
    Q => R1IN_2_1F(26),
    D => R1IN_2_1F_0(26),
    C => CLK,
    CE => EN);
\R1IN_2_1[27]\: FDE port map (
    Q => R1IN_2_1F(27),
    D => R1IN_2_1F_0(27),
    C => CLK,
    CE => EN);
\R1IN_2_1[28]\: FDE port map (
    Q => R1IN_2_1F(28),
    D => R1IN_2_1F_0(28),
    C => CLK,
    CE => EN);
\R1IN_2_1[29]\: FDE port map (
    Q => R1IN_2_1F(29),
    D => R1IN_2_1F_0(29),
    C => CLK,
    CE => EN);
\R1IN_2_1[30]\: FDE port map (
    Q => R1IN_2_1F(30),
    D => R1IN_2_1F_0(30),
    C => CLK,
    CE => EN);
\R1IN_2_1[31]\: FDE port map (
    Q => R1IN_2_1F(31),
    D => R1IN_2_1F_0(31),
    C => CLK,
    CE => EN);
\R1IN_2_1[32]\: FDE port map (
    Q => R1IN_2_1F(32),
    D => R1IN_2_1F_0(32),
    C => CLK,
    CE => EN);
\R1IN_2_1[33]\: FDE port map (
    Q => R1IN_2_1F(33),
    D => R1IN_2_1F_0(33),
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_Z5917: FDE port map (
    Q => R2_PIPE_165_RET,
    D => R1IN_ADD_1_1_S_28,
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_1_Z5918: FDE port map (
    Q => R2_PIPE_165_RET_1,
    D => R1IN_ADD_1_1_0_S_28,
    C => CLK,
    CE => EN);
R2_PIPE_165_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_19,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_164_RET_Z5920: FDE port map (
    Q => R2_PIPE_164_RET,
    D => R1IN_ADD_1_1_S_27,
    C => CLK,
    CE => EN);
R2_PIPE_164_RET_1_Z5921: FDE port map (
    Q => R2_PIPE_164_RET_1,
    D => R1IN_ADD_1_1_0_S_27,
    C => CLK,
    CE => EN);
R2_PIPE_164_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_20,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_163_RET_Z5923: FDE port map (
    Q => R2_PIPE_163_RET,
    D => R1IN_ADD_1_1_S_26,
    C => CLK,
    CE => EN);
R2_PIPE_163_RET_1_Z5924: FDE port map (
    Q => R2_PIPE_163_RET_1,
    D => R1IN_ADD_1_1_0_S_26,
    C => CLK,
    CE => EN);
R2_PIPE_163_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_21,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_162_RET_Z5926: FDE port map (
    Q => R2_PIPE_162_RET,
    D => R1IN_ADD_1_1_S_25,
    C => CLK,
    CE => EN);
R2_PIPE_162_RET_1_Z5927: FDE port map (
    Q => R2_PIPE_162_RET_1,
    D => R1IN_ADD_1_1_0_S_25,
    C => CLK,
    CE => EN);
R2_PIPE_162_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_22,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_161_RET_Z5929: FDE port map (
    Q => R2_PIPE_161_RET,
    D => R1IN_ADD_1_1_S_24,
    C => CLK,
    CE => EN);
R2_PIPE_161_RET_1_Z5930: FDE port map (
    Q => R2_PIPE_161_RET_1,
    D => R1IN_ADD_1_1_0_S_24,
    C => CLK,
    CE => EN);
R2_PIPE_161_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_23,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_160_RET_Z5932: FDE port map (
    Q => R2_PIPE_160_RET,
    D => R1IN_ADD_1_1_S_23,
    C => CLK,
    CE => EN);
R2_PIPE_160_RET_1_Z5933: FDE port map (
    Q => R2_PIPE_160_RET_1,
    D => R1IN_ADD_1_1_0_S_23,
    C => CLK,
    CE => EN);
R2_PIPE_160_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_24,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_159_RET_Z5935: FDE port map (
    Q => R2_PIPE_159_RET,
    D => R1IN_ADD_1_1_S_22,
    C => CLK,
    CE => EN);
R2_PIPE_159_RET_1_Z5936: FDE port map (
    Q => R2_PIPE_159_RET_1,
    D => R1IN_ADD_1_1_0_S_22,
    C => CLK,
    CE => EN);
R2_PIPE_159_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_25,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_158_RET_Z5938: FDE port map (
    Q => R2_PIPE_158_RET,
    D => R1IN_ADD_1_1_S_21,
    C => CLK,
    CE => EN);
R2_PIPE_158_RET_1_Z5939: FDE port map (
    Q => R2_PIPE_158_RET_1,
    D => R1IN_ADD_1_1_0_S_21,
    C => CLK,
    CE => EN);
R2_PIPE_158_RET_2: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_26,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_166_RET: FDE port map (
    Q => R1IN_ADD_1_0_CRY_31_RETO_27,
    D => R1IN_ADD_1_0_CRY_31,
    C => CLK,
    CE => EN);
R2_PIPE_166_RET_1: FDE port map (
    Q => R1IN_ADD_1_1_0_CRY_28_RETO,
    D => R1IN_ADD_1_1_0_CRY_28,
    C => CLK,
    CE => EN);
R2_PIPE_166_RET_2: FDE port map (
    Q => R1IN_ADD_1_1_CRY_28_RETO,
    D => R1IN_ADD_1_1_CRY_28,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_48_Z5944: FDE port map (
    Q => R2_PIPE_104_RET_48,
    D => N_1822_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_49_Z5945: FDE port map (
    Q => R2_PIPE_104_RET_49,
    D => N_1821_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_93_Z5946: FDE port map (
    Q => R2_PIPE_104_RET_93,
    D => N_1820_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_94_Z5947: FDE port map (
    Q => R2_PIPE_104_RET_94,
    D => N_1819_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_95_Z5948: FDE port map (
    Q => R2_PIPE_104_RET_95,
    D => N_1818_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_96_Z5949: FDE port map (
    Q => R2_PIPE_104_RET_96,
    D => N_1817_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_97_Z5950: FDE port map (
    Q => R2_PIPE_104_RET_97,
    D => N_1816_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_98_Z5951: FDE port map (
    Q => R2_PIPE_104_RET_98,
    D => N_1815_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_99_Z5952: FDE port map (
    Q => R2_PIPE_104_RET_99,
    D => N_1814_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_100_Z5953: FDE port map (
    Q => R2_PIPE_104_RET_100,
    D => N_1813_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_101_Z5954: FDE port map (
    Q => R2_PIPE_104_RET_101,
    D => N_1812_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_102_Z5955: FDE port map (
    Q => R2_PIPE_104_RET_102,
    D => N_1811_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_103_Z5956: FDE port map (
    Q => R2_PIPE_104_RET_103,
    D => N_1810_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_104_Z5957: FDE port map (
    Q => R2_PIPE_104_RET_104,
    D => N_1809_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_105_Z5958: FDE port map (
    Q => R2_PIPE_104_RET_105,
    D => N_1808_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_106_Z5959: FDE port map (
    Q => R2_PIPE_104_RET_106,
    D => N_1807_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_107_Z5960: FDE port map (
    Q => R2_PIPE_104_RET_107,
    D => N_1806_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_108_Z5961: FDE port map (
    Q => R2_PIPE_104_RET_108,
    D => N_1805_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_109_Z5962: FDE port map (
    Q => R2_PIPE_104_RET_109,
    D => N_1804_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_110_Z5963: FDE port map (
    Q => R2_PIPE_104_RET_110,
    D => N_1803_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_111_Z5964: FDE port map (
    Q => R2_PIPE_104_RET_111,
    D => N_1802_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_112_Z5965: FDE port map (
    Q => R2_PIPE_104_RET_112,
    D => N_1801_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_113_Z5966: FDE port map (
    Q => R2_PIPE_104_RET_113,
    D => N_1800_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_114_Z5967: FDE port map (
    Q => R2_PIPE_104_RET_114,
    D => N_1799_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_115_Z5968: FDE port map (
    Q => R2_PIPE_104_RET_115,
    D => N_1798_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_116_Z5969: FDE port map (
    Q => R2_PIPE_104_RET_116,
    D => N_1797_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_117_Z5970: FDE port map (
    Q => R2_PIPE_104_RET_117,
    D => N_1796_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_118_Z5971: FDE port map (
    Q => R2_PIPE_104_RET_118,
    D => N_1795_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_119_Z5972: FDE port map (
    Q => R2_PIPE_104_RET_119,
    D => N_1794_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_120_Z5973: FDE port map (
    Q => R2_PIPE_104_RET_120,
    D => N_1793_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_121_Z5974: FDE port map (
    Q => R2_PIPE_104_RET_121,
    D => N_1792_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_122_Z5975: FDE port map (
    Q => R2_PIPE_104_RET_122,
    D => N_1791_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_123_Z5976: FDE port map (
    Q => R2_PIPE_104_RET_123,
    D => N_1790_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_124_Z5977: FDE port map (
    Q => R2_PIPE_104_RET_124,
    D => N_1789_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_125: FDE port map (
    Q => R1IN_4_ADD_2_1_0_AXB_0_RETO,
    D => R1IN_4_ADD_2_1_0_AXB_0_RET_0I,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1027_Z5979: FDE port map (
    Q => R2_PIPE_104_RET_1027,
    D => N_1781_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1028_Z5980: FDE port map (
    Q => R2_PIPE_104_RET_1028,
    D => N_1779_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1029_Z5981: FDE port map (
    Q => R2_PIPE_104_RET_1029,
    D => N_1777_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1030_Z5982: FDE port map (
    Q => R2_PIPE_104_RET_1030,
    D => N_1775_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1031_Z5983: FDE port map (
    Q => R2_PIPE_104_RET_1031,
    D => N_1773_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1032_Z5984: FDE port map (
    Q => R2_PIPE_104_RET_1032,
    D => N_1771_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1033_Z5985: FDE port map (
    Q => R2_PIPE_104_RET_1033,
    D => N_1769_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1034_Z5986: FDE port map (
    Q => R2_PIPE_104_RET_1034,
    D => N_1767_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1035_Z5987: FDE port map (
    Q => R2_PIPE_104_RET_1035,
    D => N_1765_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1036_Z5988: FDE port map (
    Q => R2_PIPE_104_RET_1036,
    D => N_1763_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1037_Z5989: FDE port map (
    Q => R2_PIPE_104_RET_1037,
    D => N_1761_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1038_Z5990: FDE port map (
    Q => R2_PIPE_104_RET_1038,
    D => N_1759_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1039_Z5991: FDE port map (
    Q => R2_PIPE_104_RET_1039,
    D => N_1757_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1040_Z5992: FDE port map (
    Q => R2_PIPE_104_RET_1040,
    D => N_1755_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1041_Z5993: FDE port map (
    Q => R2_PIPE_104_RET_1041,
    D => N_1753_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1042_Z5994: FDE port map (
    Q => R2_PIPE_104_RET_1042,
    D => N_1751_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1043_Z5995: FDE port map (
    Q => R2_PIPE_104_RET_1043,
    D => N_1749_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1044_Z5996: FDE port map (
    Q => R2_PIPE_104_RET_1044,
    D => N_1747_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1045_Z5997: FDE port map (
    Q => R2_PIPE_104_RET_1045,
    D => N_1745_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1046_Z5998: FDE port map (
    Q => R2_PIPE_104_RET_1046,
    D => N_1743_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1047_Z5999: FDE port map (
    Q => R2_PIPE_104_RET_1047,
    D => N_1741_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1048_Z6000: FDE port map (
    Q => R2_PIPE_104_RET_1048,
    D => N_1739_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1049_Z6001: FDE port map (
    Q => R2_PIPE_104_RET_1049,
    D => N_1737_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1050_Z6002: FDE port map (
    Q => R2_PIPE_104_RET_1050,
    D => N_1735_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1051_Z6003: FDE port map (
    Q => R2_PIPE_104_RET_1051,
    D => N_1733_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1052_Z6004: FDE port map (
    Q => R2_PIPE_104_RET_1052,
    D => N_1731_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1053_Z6005: FDE port map (
    Q => R2_PIPE_104_RET_1053,
    D => N_1729_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1054_Z6006: FDE port map (
    Q => R2_PIPE_104_RET_1054,
    D => N_1727_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1055_Z6007: FDE port map (
    Q => R2_PIPE_104_RET_1055,
    D => N_1725_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1056_Z6008: FDE port map (
    Q => R2_PIPE_104_RET_1056,
    D => N_1723_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1057_Z6009: FDE port map (
    Q => R2_PIPE_104_RET_1057,
    D => N_1721_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1058_Z6010: FDE port map (
    Q => R2_PIPE_104_RET_1058,
    D => N_1719_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1059_Z6011: FDE port map (
    Q => R2_PIPE_104_RET_1059,
    D => N_1717_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1060_Z6012: FDE port map (
    Q => R2_PIPE_104_RET_1060,
    D => N_1715_RETI,
    C => CLK,
    CE => EN);
R2_PIPE_104_RET_1061: FDE port map (
    Q => R1IN_4_ADD_2_1_AXB_0,
    D => R1IN_4_ADD_2_1_AXB_0_RETI,
    C => CLK,
    CE => EN);
R1IN_ADD_1_1_CRY_28_Z6014: MUXCY port map (
    DI => R1IN_3(60),
    CI => R1IN_ADD_1_1_CRY_27,
    S => R1IN_ADD_1_1_AXB_28,
    O => R1IN_ADD_1_1_CRY_28);
R1IN_ADD_2_1_0_AXB_0_Z6015: LUT4 
generic map(
  INIT => X"596A"
)
port map (
  I0 => R1IN_4F(36),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_26,
  I2 => R2_PIPE_158_RET_1,
  I3 => R2_PIPE_158_RET,
  O => R1IN_ADD_2_1_0_AXB_0);
R1IN_ADD_2_1_AXB_0_Z6016: LUT4 
generic map(
  INIT => X"596A"
)
port map (
  I0 => R1IN_4F(36),
  I1 => R1IN_ADD_1_0_CRY_31_RETO_26,
  I2 => R2_PIPE_158_RET_1,
  I3 => R2_PIPE_158_RET,
  O => R1IN_ADD_2_1_AXB_0);
R1IN_ADD_2_1_AXB_51_Z6017: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO,
  I1 => R2_PIPE_104_RET_48,
  I2 => R2_PIPE_104_RET_1027,
  O => R1IN_ADD_2_1_AXB_51);
R1IN_ADD_2_1_0_AXB_51_Z6018: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => R1IN_4_ADD_2_0_CRY_35_RETO,
  I1 => R2_PIPE_104_RET_48,
  I2 => R2_PIPE_104_RET_1027,
  O => R1IN_ADD_2_1_0_AXB_51);
R1IN_4_ADD_2_1_0_S_34: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_34,
    CI => R1IN_4_ADD_2_1_0_CRY_33,
    O => N_1822_RET_0I);
R1IN_4_ADD_2_1_0_AXB_34_Z7179: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(53),
  LO => R1IN_4_ADD_2_1_0_AXB_34);
R1IN_4_ADD_2_1_0_CRY_33_Z7180: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_32,
    S => R1IN_4_ADD_2_1_0_AXB_33,
    LO => R1IN_4_ADD_2_1_0_CRY_33);
R1IN_4_ADD_2_1_0_CRY_32_Z7181: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_31,
    S => R1IN_4_ADD_2_1_0_AXB_32,
    LO => R1IN_4_ADD_2_1_0_CRY_32);
R1IN_4_ADD_2_1_0_S_33: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_33,
    CI => R1IN_4_ADD_2_1_0_CRY_32,
    O => N_1821_RET_0I);
R1IN_4_ADD_2_1_0_AXB_33_Z7183: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(52),
  LO => R1IN_4_ADD_2_1_0_AXB_33);
R1IN_4_ADD_2_1_0_CRY_31_Z7184: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_30,
    S => R1IN_4_ADD_2_1_0_AXB_31,
    LO => R1IN_4_ADD_2_1_0_CRY_31);
R1IN_4_ADD_2_1_0_S_32: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_32,
    CI => R1IN_4_ADD_2_1_0_CRY_31,
    O => N_1820_RET_0I);
R1IN_4_ADD_2_1_0_AXB_32_Z7186: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(51),
  LO => R1IN_4_ADD_2_1_0_AXB_32);
R1IN_4_ADD_2_1_0_CRY_30_Z7187: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_29,
    S => R1IN_4_ADD_2_1_0_AXB_30,
    LO => R1IN_4_ADD_2_1_0_CRY_30);
R1IN_4_ADD_2_1_0_S_31: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_31,
    CI => R1IN_4_ADD_2_1_0_CRY_30,
    O => N_1819_RET_0I);
R1IN_4_ADD_2_1_0_AXB_31_Z7189: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(50),
  LO => R1IN_4_ADD_2_1_0_AXB_31);
R1IN_4_ADD_2_1_0_CRY_29_Z7190: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_28,
    S => R1IN_4_ADD_2_1_0_AXB_29,
    LO => R1IN_4_ADD_2_1_0_CRY_29);
R1IN_4_ADD_2_1_0_S_30: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_30,
    CI => R1IN_4_ADD_2_1_0_CRY_29,
    O => N_1818_RET_0I);
R1IN_4_ADD_2_1_0_AXB_30_Z7192: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(49),
  LO => R1IN_4_ADD_2_1_0_AXB_30);
R1IN_4_ADD_2_1_0_CRY_28_Z7193: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_27,
    S => R1IN_4_ADD_2_1_0_AXB_28,
    LO => R1IN_4_ADD_2_1_0_CRY_28);
R1IN_4_ADD_2_1_0_S_29: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_29,
    CI => R1IN_4_ADD_2_1_0_CRY_28,
    O => N_1817_RET_0I);
R1IN_4_ADD_2_1_0_AXB_29_Z7195: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(48),
  LO => R1IN_4_ADD_2_1_0_AXB_29);
R1IN_4_ADD_2_1_0_CRY_27_Z7196: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_26,
    S => R1IN_4_ADD_2_1_0_AXB_27,
    LO => R1IN_4_ADD_2_1_0_CRY_27);
R1IN_4_ADD_2_1_0_S_28: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_28,
    CI => R1IN_4_ADD_2_1_0_CRY_27,
    O => N_1816_RET_0I);
R1IN_4_ADD_2_1_0_AXB_28_Z7198: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(47),
  LO => R1IN_4_ADD_2_1_0_AXB_28);
R1IN_4_ADD_2_1_0_CRY_26_Z7199: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_25,
    S => R1IN_4_ADD_2_1_0_AXB_26,
    LO => R1IN_4_ADD_2_1_0_CRY_26);
R1IN_4_ADD_2_1_0_S_27: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_27,
    CI => R1IN_4_ADD_2_1_0_CRY_26,
    O => N_1815_RET_0I);
R1IN_4_ADD_2_1_0_AXB_27_Z7201: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(46),
  LO => R1IN_4_ADD_2_1_0_AXB_27);
R1IN_4_ADD_2_1_0_CRY_25_Z7202: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_24,
    S => R1IN_4_ADD_2_1_0_AXB_25,
    LO => R1IN_4_ADD_2_1_0_CRY_25);
R1IN_4_ADD_2_1_0_S_26: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_26,
    CI => R1IN_4_ADD_2_1_0_CRY_25,
    O => N_1814_RET_0I);
R1IN_4_ADD_2_1_0_AXB_26_Z7204: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(45),
  LO => R1IN_4_ADD_2_1_0_AXB_26);
R1IN_4_ADD_2_1_0_CRY_24_Z7205: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_23,
    S => R1IN_4_ADD_2_1_0_AXB_24,
    LO => R1IN_4_ADD_2_1_0_CRY_24);
R1IN_4_ADD_2_1_0_S_25: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_25,
    CI => R1IN_4_ADD_2_1_0_CRY_24,
    O => N_1813_RET_0I);
R1IN_4_ADD_2_1_0_AXB_25_Z7207: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(44),
  LO => R1IN_4_ADD_2_1_0_AXB_25);
R1IN_4_ADD_2_1_0_CRY_23_Z7208: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_22,
    S => R1IN_4_ADD_2_1_0_AXB_23,
    LO => R1IN_4_ADD_2_1_0_CRY_23);
R1IN_4_ADD_2_1_0_S_24: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_24,
    CI => R1IN_4_ADD_2_1_0_CRY_23,
    O => N_1812_RET_0I);
R1IN_4_ADD_2_1_0_AXB_24_Z7210: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(43),
  LO => R1IN_4_ADD_2_1_0_AXB_24);
R1IN_4_ADD_2_1_0_CRY_22_Z7211: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_21,
    S => R1IN_4_ADD_2_1_0_AXB_22,
    LO => R1IN_4_ADD_2_1_0_CRY_22);
R1IN_4_ADD_2_1_0_S_23: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_23,
    CI => R1IN_4_ADD_2_1_0_CRY_22,
    O => N_1811_RET_0I);
R1IN_4_ADD_2_1_0_AXB_23_Z7213: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(42),
  LO => R1IN_4_ADD_2_1_0_AXB_23);
R1IN_4_ADD_2_1_0_CRY_21_Z7214: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_20,
    S => R1IN_4_ADD_2_1_0_AXB_21,
    LO => R1IN_4_ADD_2_1_0_CRY_21);
R1IN_4_ADD_2_1_0_S_22: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_22,
    CI => R1IN_4_ADD_2_1_0_CRY_21,
    O => N_1810_RET_0I);
R1IN_4_ADD_2_1_0_AXB_22_Z7216: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(41),
  LO => R1IN_4_ADD_2_1_0_AXB_22);
R1IN_4_ADD_2_1_0_CRY_20_Z7217: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_19,
    S => R1IN_4_ADD_2_1_0_AXB_20,
    LO => R1IN_4_ADD_2_1_0_CRY_20);
R1IN_4_ADD_2_1_0_S_21: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_21,
    CI => R1IN_4_ADD_2_1_0_CRY_20,
    O => N_1809_RET_0I);
R1IN_4_ADD_2_1_0_AXB_21_Z7219: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(40),
  LO => R1IN_4_ADD_2_1_0_AXB_21);
R1IN_4_ADD_2_1_0_CRY_19_Z7220: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_18,
    S => R1IN_4_ADD_2_1_0_AXB_19,
    LO => R1IN_4_ADD_2_1_0_CRY_19);
R1IN_4_ADD_2_1_0_S_20: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_20,
    CI => R1IN_4_ADD_2_1_0_CRY_19,
    O => N_1808_RET_0I);
R1IN_4_ADD_2_1_0_AXB_20_Z7222: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(39),
  LO => R1IN_4_ADD_2_1_0_AXB_20);
R1IN_4_ADD_2_1_0_CRY_18_Z7223: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_17,
    S => R1IN_4_ADD_2_1_0_AXB_18,
    LO => R1IN_4_ADD_2_1_0_CRY_18);
R1IN_4_ADD_2_1_0_S_19: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_19,
    CI => R1IN_4_ADD_2_1_0_CRY_18,
    O => N_1807_RET_0I);
R1IN_4_ADD_2_1_0_AXB_19_Z7225: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(38),
  LO => R1IN_4_ADD_2_1_0_AXB_19);
R1IN_4_ADD_2_1_0_CRY_17_Z7226: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_16,
    S => R1IN_4_ADD_2_1_0_AXB_17,
    LO => R1IN_4_ADD_2_1_0_CRY_17);
R1IN_4_ADD_2_1_0_S_18: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_18,
    CI => R1IN_4_ADD_2_1_0_CRY_17,
    O => N_1806_RET_0I);
R1IN_4_ADD_2_1_0_AXB_18_Z7228: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(37),
  LO => R1IN_4_ADD_2_1_0_AXB_18);
R1IN_4_ADD_2_1_0_CRY_16_Z7229: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_15,
    S => R1IN_4_ADD_2_1_0_AXB_16,
    LO => R1IN_4_ADD_2_1_0_CRY_16);
R1IN_4_ADD_2_1_0_S_17: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_17,
    CI => R1IN_4_ADD_2_1_0_CRY_16,
    O => N_1805_RET_0I);
R1IN_4_ADD_2_1_0_AXB_17_Z7231: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(36),
  LO => R1IN_4_ADD_2_1_0_AXB_17);
R1IN_4_ADD_2_1_0_CRY_15_Z7232: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_14,
    S => R1IN_4_ADD_2_1_0_AXB_15,
    LO => R1IN_4_ADD_2_1_0_CRY_15);
R1IN_4_ADD_2_1_0_S_16: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_16,
    CI => R1IN_4_ADD_2_1_0_CRY_15,
    O => N_1804_RET_0I);
R1IN_4_ADD_2_1_0_AXB_16_Z7234: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(35),
  LO => R1IN_4_ADD_2_1_0_AXB_16);
R1IN_4_ADD_2_1_0_CRY_14_Z7235: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_13,
    S => R1IN_4_ADD_2_1_0_AXB_14,
    LO => R1IN_4_ADD_2_1_0_CRY_14);
R1IN_4_ADD_2_1_0_S_15: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_15,
    CI => R1IN_4_ADD_2_1_0_CRY_14,
    O => N_1803_RET_0I);
R1IN_4_ADD_2_1_0_AXB_15_Z7237: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(34),
  LO => R1IN_4_ADD_2_1_0_AXB_15);
R1IN_4_ADD_2_1_0_CRY_13_Z7238: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_12,
    S => R1IN_4_ADD_2_1_0_AXB_13,
    LO => R1IN_4_ADD_2_1_0_CRY_13);
R1IN_4_ADD_2_1_0_S_14: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_14,
    CI => R1IN_4_ADD_2_1_0_CRY_13,
    O => N_1802_RET_0I);
R1IN_4_ADD_2_1_0_AXB_14_Z7240: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(33),
  LO => R1IN_4_ADD_2_1_0_AXB_14);
R1IN_4_ADD_2_1_0_CRY_12_Z7241: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_11,
    S => R1IN_4_ADD_2_1_0_AXB_12,
    LO => R1IN_4_ADD_2_1_0_CRY_12);
R1IN_4_ADD_2_1_0_S_13: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_13,
    CI => R1IN_4_ADD_2_1_0_CRY_12,
    O => N_1801_RET_0I);
R1IN_4_ADD_2_1_0_AXB_13_Z7243: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(32),
  LO => R1IN_4_ADD_2_1_0_AXB_13);
R1IN_4_ADD_2_1_0_CRY_11_Z7244: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_10,
    S => R1IN_4_ADD_2_1_0_AXB_11,
    LO => R1IN_4_ADD_2_1_0_CRY_11);
R1IN_4_ADD_2_1_0_S_12: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_12,
    CI => R1IN_4_ADD_2_1_0_CRY_11,
    O => N_1800_RET_0I);
R1IN_4_ADD_2_1_0_AXB_12_Z7246: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(31),
  LO => R1IN_4_ADD_2_1_0_AXB_12);
R1IN_4_ADD_2_1_0_CRY_10_Z7247: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_9,
    S => R1IN_4_ADD_2_1_0_AXB_10,
    LO => R1IN_4_ADD_2_1_0_CRY_10);
R1IN_4_ADD_2_1_0_S_11: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_11,
    CI => R1IN_4_ADD_2_1_0_CRY_10,
    O => N_1799_RET_0I);
R1IN_4_ADD_2_1_0_AXB_11_Z7249: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(30),
  LO => R1IN_4_ADD_2_1_0_AXB_11);
R1IN_4_ADD_2_1_0_CRY_9_Z7250: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_0_CRY_8,
    S => R1IN_4_ADD_2_1_0_AXB_9,
    LO => R1IN_4_ADD_2_1_0_CRY_9);
R1IN_4_ADD_2_1_0_S_10: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_10,
    CI => R1IN_4_ADD_2_1_0_CRY_9,
    O => N_1798_RET_0I);
R1IN_4_ADD_2_1_0_AXB_10_Z7252: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(29),
  LO => R1IN_4_ADD_2_1_0_AXB_10);
R1IN_4_ADD_2_1_0_CRY_8_Z7253: MUXCY_L port map (
    DI => NN_10,
    CI => R1IN_4_ADD_2_1_0_CRY_7,
    S => R1IN_4_ADD_2_1_0_AXB_8,
    LO => R1IN_4_ADD_2_1_0_CRY_8);
R1IN_4_ADD_2_1_0_S_9: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_9,
    CI => R1IN_4_ADD_2_1_0_CRY_8,
    O => N_1797_RET_0I);
R1IN_4_ADD_2_1_0_AXB_9_Z7255: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(28),
  LO => R1IN_4_ADD_2_1_0_AXB_9);
R1IN_4_ADD_2_1_0_CRY_7_Z7256: MUXCY_L port map (
    DI => NN_9,
    CI => R1IN_4_ADD_2_1_0_CRY_6,
    S => R1IN_4_ADD_2_1_0_AXB_7,
    LO => R1IN_4_ADD_2_1_0_CRY_7);
R1IN_4_ADD_2_1_0_S_8: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_8,
    CI => R1IN_4_ADD_2_1_0_CRY_7,
    O => N_1796_RET_0I);
R1IN_4_ADD_2_1_0_AXB_8_Z7258: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(27),
  I1 => NN_10,
  LO => R1IN_4_ADD_2_1_0_AXB_8);
R1IN_4_ADD_2_1_0_CRY_6_Z7259: MUXCY_L port map (
    DI => NN_8,
    CI => R1IN_4_ADD_2_1_0_CRY_5,
    S => R1IN_4_ADD_2_1_0_AXB_6,
    LO => R1IN_4_ADD_2_1_0_CRY_6);
R1IN_4_ADD_2_1_0_S_7: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_7,
    CI => R1IN_4_ADD_2_1_0_CRY_6,
    O => N_1795_RET_0I);
R1IN_4_ADD_2_1_0_AXB_7_Z7261: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(26),
  I1 => NN_9,
  LO => R1IN_4_ADD_2_1_0_AXB_7);
R1IN_4_ADD_2_1_0_CRY_5_Z7262: MUXCY_L port map (
    DI => NN_7,
    CI => R1IN_4_ADD_2_1_0_CRY_4,
    S => R1IN_4_ADD_2_1_0_AXB_5,
    LO => R1IN_4_ADD_2_1_0_CRY_5);
R1IN_4_ADD_2_1_0_S_6: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_6,
    CI => R1IN_4_ADD_2_1_0_CRY_5,
    O => N_1794_RET_0I);
R1IN_4_ADD_2_1_0_AXB_6_Z7264: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(25),
  I1 => NN_8,
  LO => R1IN_4_ADD_2_1_0_AXB_6);
R1IN_4_ADD_2_1_0_CRY_4_Z7265: MUXCY_L port map (
    DI => NN_6,
    CI => R1IN_4_ADD_2_1_0_CRY_3,
    S => R1IN_4_ADD_2_1_0_AXB_4,
    LO => R1IN_4_ADD_2_1_0_CRY_4);
R1IN_4_ADD_2_1_0_S_5: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_5,
    CI => R1IN_4_ADD_2_1_0_CRY_4,
    O => N_1793_RET_0I);
R1IN_4_ADD_2_1_0_AXB_5_Z7267: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(24),
  I1 => NN_7,
  LO => R1IN_4_ADD_2_1_0_AXB_5);
R1IN_4_ADD_2_1_0_CRY_3_Z7268: MUXCY_L port map (
    DI => NN_5,
    CI => R1IN_4_ADD_2_1_0_CRY_2,
    S => R1IN_4_ADD_2_1_0_AXB_3,
    LO => R1IN_4_ADD_2_1_0_CRY_3);
R1IN_4_ADD_2_1_0_S_4: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_4,
    CI => R1IN_4_ADD_2_1_0_CRY_3,
    O => N_1792_RET_0I);
R1IN_4_ADD_2_1_0_AXB_4_Z7270: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(23),
  I1 => NN_6,
  LO => R1IN_4_ADD_2_1_0_AXB_4);
R1IN_4_ADD_2_1_0_CRY_2_Z7271: MUXCY_L port map (
    DI => NN_4,
    CI => R1IN_4_ADD_2_1_0_CRY_1,
    S => R1IN_4_ADD_2_1_0_AXB_2,
    LO => R1IN_4_ADD_2_1_0_CRY_2);
R1IN_4_ADD_2_1_0_S_3: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_3,
    CI => R1IN_4_ADD_2_1_0_CRY_2,
    O => N_1791_RET_0I);
R1IN_4_ADD_2_1_0_AXB_3_Z7273: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(22),
  I1 => NN_5,
  LO => R1IN_4_ADD_2_1_0_AXB_3);
R1IN_4_ADD_2_1_0_CRY_1_Z7274: MUXCY_L port map (
    DI => NN_3,
    CI => R1IN_4_ADD_2_1_0_CRY_0,
    S => R1IN_4_ADD_2_1_0_AXB_1,
    LO => R1IN_4_ADD_2_1_0_CRY_1);
R1IN_4_ADD_2_1_0_S_2: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_2,
    CI => R1IN_4_ADD_2_1_0_CRY_1,
    O => N_1790_RET_0I);
R1IN_4_ADD_2_1_0_AXB_2_Z7276: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(21),
  I1 => NN_4,
  LO => R1IN_4_ADD_2_1_0_AXB_2);
R1IN_4_ADD_2_1_0_CRY_0_Z7277: MUXCY_L port map (
    DI => R1IN_4_ADD_2_1,
    CI => NN_2,
    S => R1IN_4_ADD_2_1_0_AXB_0_RET_0I,
    LO => R1IN_4_ADD_2_1_0_CRY_0);
R1IN_4_ADD_2_1_0_S_1: XORCY port map (
    LI => R1IN_4_ADD_2_1_0_AXB_1,
    CI => R1IN_4_ADD_2_1_0_CRY_0,
    O => N_1789_RET_0I);
R1IN_4_ADD_2_1_0_AXB_1_Z7279: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(20),
  I1 => NN_3,
  LO => R1IN_4_ADD_2_1_0_AXB_1);
R1IN_4_ADD_2_1_0_AXB_0: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(19),
  I1 => R1IN_4_ADD_2_1,
  O => R1IN_4_ADD_2_1_0_AXB_0_RET_0I);
\R1IN_ADD_2_MUX[0]\: LUT3 
generic map(
  INIT => X"72"
)
port map (
  I0 => R1IN_ADD_2_0_CRY_52,
  I1 => R1IN_ADD_2_1_0_AXB_0,
  I2 => R1IN_ADD_2_1_AXB_0,
  O => PRODUCT(70));
\R1IN_ADD_1_MUX[0]\: LUT3_L 
generic map(
  INIT => X"72"
)
port map (
  I0 => R1IN_ADD_1_0_CRY_31,
  I1 => R1IN_ADD_1_1_0_AXB_0,
  I2 => R1IN_ADD_1_1_AXB_0,
  LO => R1IN_ADD_1(32));
R1IN_ADD_1_0_AXB_17_Z7371: LUT4_L 
generic map(
  INIT => X"6996"
)
port map (
  I0 => R1IN_2_1F(17),
  I1 => R1IN_2_ADD_1,
  I2 => R1IN_3_1F(17),
  I3 => R1IN_3_ADD_1,
  LO => R1IN_ADD_1_0_AXB_17);
R1IN_4_ADD_2_0_AXB_34_Z7372: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(17),
  I1 => R1IN_4_ADD_1(34),
  LO => R1IN_4_ADD_2_0_AXB_34);
\R1IN_4_ADD_2_MUX[1]\: LUT3_L 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R2_PIPE_104_RET_1060,
  I1 => R2_PIPE_104_RET_124,
  I2 => R1IN_4_ADD_2_0_CRY_35_RETO_32,
  LO => R1IN_4(54));
\R1IN_ADD_2_MUX[51]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_51,
  I1 => R1IN_ADD_2_1_0_S_51,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(121));
\R1IN_ADD_2_MUX[50]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_50,
  I1 => R1IN_ADD_2_1_0_S_50,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(120));
\R1IN_ADD_2_MUX[49]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_49,
  I1 => R1IN_ADD_2_1_0_S_49,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(119));
\R1IN_ADD_2_MUX[48]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_48,
  I1 => R1IN_ADD_2_1_0_S_48,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(118));
\R1IN_ADD_2_MUX[47]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_47,
  I1 => R1IN_ADD_2_1_0_S_47,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(117));
\R1IN_ADD_2_MUX[46]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_46,
  I1 => R1IN_ADD_2_1_0_S_46,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(116));
\R1IN_ADD_2_MUX[45]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_45,
  I1 => R1IN_ADD_2_1_0_S_45,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(115));
\R1IN_ADD_2_MUX[44]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_44,
  I1 => R1IN_ADD_2_1_0_S_44,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(114));
\R1IN_ADD_2_MUX[43]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_43,
  I1 => R1IN_ADD_2_1_0_S_43,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(113));
\R1IN_ADD_2_MUX[42]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_42,
  I1 => R1IN_ADD_2_1_0_S_42,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(112));
\R1IN_ADD_2_MUX[41]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_41,
  I1 => R1IN_ADD_2_1_0_S_41,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(111));
\R1IN_ADD_2_MUX[40]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_40,
  I1 => R1IN_ADD_2_1_0_S_40,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(110));
\R1IN_ADD_2_MUX[39]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_39,
  I1 => R1IN_ADD_2_1_0_S_39,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(109));
\R1IN_ADD_2_MUX[38]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_38,
  I1 => R1IN_ADD_2_1_0_S_38,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(108));
\R1IN_ADD_2_MUX[37]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_37,
  I1 => R1IN_ADD_2_1_0_S_37,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(107));
\R1IN_ADD_2_MUX[36]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_36,
  I1 => R1IN_ADD_2_1_0_S_36,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(106));
\R1IN_ADD_2_MUX[35]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_35,
  I1 => R1IN_ADD_2_1_0_S_35,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(105));
\R1IN_ADD_2_MUX[34]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_34,
  I1 => R1IN_ADD_2_1_0_S_34,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(104));
\R1IN_ADD_2_MUX[33]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_33,
  I1 => R1IN_ADD_2_1_0_S_33,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(103));
\R1IN_ADD_2_MUX[32]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_32,
  I1 => R1IN_ADD_2_1_0_S_32,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(102));
\R1IN_ADD_2_MUX[31]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_31,
  I1 => R1IN_ADD_2_1_0_S_31,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(101));
\R1IN_ADD_2_MUX[30]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_30,
  I1 => R1IN_ADD_2_1_0_S_30,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(100));
\R1IN_ADD_2_MUX[29]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_29,
  I1 => R1IN_ADD_2_1_0_S_29,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(99));
\R1IN_ADD_2_MUX[28]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_28,
  I1 => R1IN_ADD_2_1_0_S_28,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(98));
\R1IN_ADD_2_MUX[27]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_27,
  I1 => R1IN_ADD_2_1_0_S_27,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(97));
\R1IN_ADD_2_MUX[26]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_26,
  I1 => R1IN_ADD_2_1_0_S_26,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(96));
\R1IN_ADD_2_MUX[25]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_25,
  I1 => R1IN_ADD_2_1_0_S_25,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(95));
\R1IN_ADD_2_MUX[24]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_24,
  I1 => R1IN_ADD_2_1_0_S_24,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(94));
\R1IN_ADD_2_MUX[23]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_23,
  I1 => R1IN_ADD_2_1_0_S_23,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(93));
\R1IN_ADD_2_MUX[22]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_22,
  I1 => R1IN_ADD_2_1_0_S_22,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(92));
\R1IN_ADD_2_MUX[21]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_21,
  I1 => R1IN_ADD_2_1_0_S_21,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(91));
\R1IN_ADD_2_MUX[20]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_20,
  I1 => R1IN_ADD_2_1_0_S_20,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(90));
\R1IN_ADD_2_MUX[19]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_19,
  I1 => R1IN_ADD_2_1_0_S_19,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(89));
\R1IN_ADD_2_MUX[18]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_18,
  I1 => R1IN_ADD_2_1_0_S_18,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(88));
\R1IN_ADD_2_MUX[17]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_17,
  I1 => R1IN_ADD_2_1_0_S_17,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(87));
\R1IN_ADD_2_MUX[16]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_16,
  I1 => R1IN_ADD_2_1_0_S_16,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(86));
\R1IN_ADD_2_MUX[15]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_15,
  I1 => R1IN_ADD_2_1_0_S_15,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(85));
\R1IN_ADD_2_MUX[14]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_14,
  I1 => R1IN_ADD_2_1_0_S_14,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(84));
\R1IN_ADD_2_MUX[13]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_13,
  I1 => R1IN_ADD_2_1_0_S_13,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(83));
\R1IN_ADD_2_MUX[12]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_12,
  I1 => R1IN_ADD_2_1_0_S_12,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(82));
\R1IN_ADD_2_MUX[11]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_11,
  I1 => R1IN_ADD_2_1_0_S_11,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(81));
\R1IN_ADD_2_MUX[10]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_10,
  I1 => R1IN_ADD_2_1_0_S_10,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(80));
\R1IN_ADD_2_MUX[9]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_9,
  I1 => R1IN_ADD_2_1_0_S_9,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(79));
\R1IN_ADD_2_MUX[8]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_8,
  I1 => R1IN_ADD_2_1_0_S_8,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(78));
\R1IN_ADD_2_MUX[7]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_7,
  I1 => R1IN_ADD_2_1_0_S_7,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(77));
\R1IN_ADD_2_MUX[6]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_6,
  I1 => R1IN_ADD_2_1_0_S_6,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(76));
\R1IN_ADD_2_MUX[5]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_5,
  I1 => R1IN_ADD_2_1_0_S_5,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(75));
\R1IN_ADD_2_MUX[4]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_4,
  I1 => R1IN_ADD_2_1_0_S_4,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(74));
\R1IN_ADD_2_MUX[3]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_3,
  I1 => R1IN_ADD_2_1_0_S_3,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(73));
\R1IN_ADD_2_MUX[2]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_2,
  I1 => R1IN_ADD_2_1_0_S_2,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(72));
\R1IN_ADD_2_MUX[1]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => R1IN_ADD_2_1_S_1,
  I1 => R1IN_ADD_2_1_0_S_1,
  I2 => R1IN_ADD_2_0_CRY_52,
  O => PRODUCT(71));
R1IN_4_ADD_1_AXB_0: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_3F(0),
  I1 => NN_12,
  O => R1IN_4_ADD_2_0);
R1IN_4_4_ADD_2_AXB_36_Z7426: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4_4F(19),
  O => R1IN_4_4_ADD_2_AXB_36);
R1IN_4_4_ADD_2_AXB_0: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4_ADD_1F(0),
  I1 => R1IN_4_4_ADD_2,
  O => R1IN_4_4(17));
R1IN_2_ADD_1_AXB_43_Z7428: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_2_2F(43),
  O => R1IN_2_ADD_1_AXB_43);
R1IN_3_ADD_1_AXB_43_Z7429: LUT1 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_3_2F(43),
  O => R1IN_3_ADD_1_AXB_43);
R1IN_3_ADD_1_AXB_0: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_3_1F(17),
  I1 => R1IN_3_ADD_1,
  O => R1IN_3(17));
R1IN_ADD_1_1_0_AXB_28_Z7431: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(60),
  I1 => R1IN_3(60),
  LO => R1IN_ADD_1_1_0_AXB_28);
R1IN_ADD_1_1_0_AXB_27_Z7432: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(59),
  I1 => R1IN_3(59),
  LO => R1IN_ADD_1_1_0_AXB_27);
R1IN_ADD_1_1_0_AXB_26_Z7433: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(58),
  I1 => R1IN_3(58),
  LO => R1IN_ADD_1_1_0_AXB_26);
R1IN_ADD_1_1_0_AXB_25_Z7434: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(57),
  I1 => R1IN_3(57),
  LO => R1IN_ADD_1_1_0_AXB_25);
R1IN_ADD_1_1_0_AXB_24_Z7435: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(56),
  I1 => R1IN_3(56),
  LO => R1IN_ADD_1_1_0_AXB_24);
R1IN_ADD_1_1_0_AXB_23_Z7436: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(55),
  I1 => R1IN_3(55),
  LO => R1IN_ADD_1_1_0_AXB_23);
R1IN_ADD_1_1_0_AXB_22_Z7437: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(54),
  I1 => R1IN_3(54),
  LO => R1IN_ADD_1_1_0_AXB_22);
R1IN_ADD_1_1_0_AXB_21_Z7438: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(53),
  I1 => R1IN_3(53),
  LO => R1IN_ADD_1_1_0_AXB_21);
R1IN_ADD_1_1_0_AXB_20_Z7439: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(52),
  I1 => R1IN_3(52),
  LO => R1IN_ADD_1_1_0_AXB_20);
R1IN_ADD_1_1_0_AXB_19_Z7440: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(51),
  I1 => R1IN_3(51),
  LO => R1IN_ADD_1_1_0_AXB_19);
R1IN_ADD_1_1_0_AXB_18_Z7441: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(50),
  I1 => R1IN_3(50),
  LO => R1IN_ADD_1_1_0_AXB_18);
R1IN_ADD_1_1_0_AXB_17_Z7442: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(49),
  I1 => R1IN_3(49),
  LO => R1IN_ADD_1_1_0_AXB_17);
R1IN_ADD_1_1_0_AXB_16_Z7443: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(48),
  I1 => R1IN_3(48),
  LO => R1IN_ADD_1_1_0_AXB_16);
R1IN_ADD_1_1_0_AXB_15_Z7444: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(47),
  I1 => R1IN_3(47),
  LO => R1IN_ADD_1_1_0_AXB_15);
R1IN_ADD_1_1_0_AXB_14_Z7445: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(46),
  I1 => R1IN_3(46),
  LO => R1IN_ADD_1_1_0_AXB_14);
R1IN_ADD_1_1_0_AXB_13_Z7446: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(45),
  I1 => R1IN_3(45),
  LO => R1IN_ADD_1_1_0_AXB_13);
R1IN_ADD_1_1_0_AXB_12_Z7447: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(44),
  I1 => R1IN_3(44),
  LO => R1IN_ADD_1_1_0_AXB_12);
R1IN_ADD_1_1_0_AXB_11_Z7448: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(43),
  I1 => R1IN_3(43),
  LO => R1IN_ADD_1_1_0_AXB_11);
R1IN_ADD_1_1_0_AXB_10_Z7449: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(42),
  I1 => R1IN_3(42),
  LO => R1IN_ADD_1_1_0_AXB_10);
R1IN_ADD_1_1_0_AXB_9_Z7450: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(41),
  I1 => R1IN_3(41),
  LO => R1IN_ADD_1_1_0_AXB_9);
R1IN_ADD_1_1_0_AXB_8_Z7451: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(40),
  I1 => R1IN_3(40),
  LO => R1IN_ADD_1_1_0_AXB_8);
R1IN_ADD_1_1_0_AXB_7_Z7452: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(39),
  I1 => R1IN_3(39),
  LO => R1IN_ADD_1_1_0_AXB_7);
R1IN_ADD_1_1_0_AXB_6_Z7453: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(38),
  I1 => R1IN_3(38),
  LO => R1IN_ADD_1_1_0_AXB_6);
R1IN_ADD_1_1_0_AXB_5_Z7454: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(37),
  I1 => R1IN_3(37),
  LO => R1IN_ADD_1_1_0_AXB_5);
R1IN_ADD_1_1_0_AXB_4_Z7455: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(36),
  I1 => R1IN_3(36),
  LO => R1IN_ADD_1_1_0_AXB_4);
R1IN_ADD_1_1_0_AXB_3_Z7456: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(35),
  I1 => R1IN_3(35),
  LO => R1IN_ADD_1_1_0_AXB_3);
R1IN_ADD_1_1_0_AXB_2_Z7457: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(34),
  I1 => R1IN_3(34),
  LO => R1IN_ADD_1_1_0_AXB_2);
R1IN_ADD_1_1_0_AXB_1_Z7458: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(33),
  I1 => R1IN_3(33),
  LO => R1IN_ADD_1_1_0_AXB_1);
R1IN_ADD_1_1_0_AXB_0_Z7459: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(32),
  I1 => R1IN_3(32),
  O => R1IN_ADD_1_1_0_AXB_0);
R1IN_ADD_1_1_AXB_28_Z7460: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(60),
  I1 => R1IN_3(60),
  LO => R1IN_ADD_1_1_AXB_28);
R1IN_ADD_1_1_AXB_27_Z7461: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(59),
  I1 => R1IN_3(59),
  LO => R1IN_ADD_1_1_AXB_27);
R1IN_ADD_1_1_AXB_26_Z7462: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(58),
  I1 => R1IN_3(58),
  LO => R1IN_ADD_1_1_AXB_26);
R1IN_ADD_1_1_AXB_25_Z7463: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(57),
  I1 => R1IN_3(57),
  LO => R1IN_ADD_1_1_AXB_25);
R1IN_ADD_1_1_AXB_24_Z7464: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(56),
  I1 => R1IN_3(56),
  LO => R1IN_ADD_1_1_AXB_24);
R1IN_ADD_1_1_AXB_23_Z7465: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(55),
  I1 => R1IN_3(55),
  LO => R1IN_ADD_1_1_AXB_23);
R1IN_ADD_1_1_AXB_22_Z7466: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(54),
  I1 => R1IN_3(54),
  LO => R1IN_ADD_1_1_AXB_22);
R1IN_ADD_1_1_AXB_21_Z7467: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(53),
  I1 => R1IN_3(53),
  LO => R1IN_ADD_1_1_AXB_21);
R1IN_ADD_1_1_AXB_20_Z7468: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(52),
  I1 => R1IN_3(52),
  LO => R1IN_ADD_1_1_AXB_20);
R1IN_ADD_1_1_AXB_19_Z7469: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(51),
  I1 => R1IN_3(51),
  LO => R1IN_ADD_1_1_AXB_19);
R1IN_ADD_1_1_AXB_18_Z7470: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(50),
  I1 => R1IN_3(50),
  LO => R1IN_ADD_1_1_AXB_18);
R1IN_ADD_1_1_AXB_17_Z7471: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(49),
  I1 => R1IN_3(49),
  LO => R1IN_ADD_1_1_AXB_17);
R1IN_ADD_1_1_AXB_16_Z7472: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(48),
  I1 => R1IN_3(48),
  LO => R1IN_ADD_1_1_AXB_16);
R1IN_ADD_1_1_AXB_15_Z7473: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(47),
  I1 => R1IN_3(47),
  LO => R1IN_ADD_1_1_AXB_15);
R1IN_ADD_1_1_AXB_14_Z7474: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(46),
  I1 => R1IN_3(46),
  LO => R1IN_ADD_1_1_AXB_14);
R1IN_ADD_1_1_AXB_13_Z7475: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(45),
  I1 => R1IN_3(45),
  LO => R1IN_ADD_1_1_AXB_13);
R1IN_ADD_1_1_AXB_12_Z7476: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(44),
  I1 => R1IN_3(44),
  LO => R1IN_ADD_1_1_AXB_12);
R1IN_ADD_1_1_AXB_11_Z7477: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(43),
  I1 => R1IN_3(43),
  LO => R1IN_ADD_1_1_AXB_11);
R1IN_ADD_1_1_AXB_10_Z7478: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(42),
  I1 => R1IN_3(42),
  LO => R1IN_ADD_1_1_AXB_10);
R1IN_ADD_1_1_AXB_9_Z7479: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(41),
  I1 => R1IN_3(41),
  LO => R1IN_ADD_1_1_AXB_9);
R1IN_ADD_1_1_AXB_8_Z7480: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(40),
  I1 => R1IN_3(40),
  LO => R1IN_ADD_1_1_AXB_8);
R1IN_ADD_1_1_AXB_7_Z7481: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(39),
  I1 => R1IN_3(39),
  LO => R1IN_ADD_1_1_AXB_7);
R1IN_ADD_1_1_AXB_6_Z7482: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(38),
  I1 => R1IN_3(38),
  LO => R1IN_ADD_1_1_AXB_6);
R1IN_ADD_1_1_AXB_5_Z7483: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(37),
  I1 => R1IN_3(37),
  LO => R1IN_ADD_1_1_AXB_5);
R1IN_ADD_1_1_AXB_4_Z7484: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(36),
  I1 => R1IN_3(36),
  LO => R1IN_ADD_1_1_AXB_4);
R1IN_ADD_1_1_AXB_3_Z7485: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(35),
  I1 => R1IN_3(35),
  LO => R1IN_ADD_1_1_AXB_3);
R1IN_ADD_1_1_AXB_2_Z7486: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(34),
  I1 => R1IN_3(34),
  LO => R1IN_ADD_1_1_AXB_2);
R1IN_ADD_1_1_AXB_1_Z7487: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(33),
  I1 => R1IN_3(33),
  LO => R1IN_ADD_1_1_AXB_1);
R1IN_ADD_1_1_AXB_0_Z7488: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(32),
  I1 => R1IN_3(32),
  O => R1IN_ADD_1_1_AXB_0);
R1IN_ADD_1_0_AXB_31_Z7489: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(31),
  I1 => R1IN_3(31),
  LO => R1IN_ADD_1_0_AXB_31);
R1IN_ADD_1_0_AXB_30_Z7490: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(30),
  I1 => R1IN_3(30),
  LO => R1IN_ADD_1_0_AXB_30);
R1IN_ADD_1_0_AXB_29_Z7491: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(29),
  I1 => R1IN_3(29),
  LO => R1IN_ADD_1_0_AXB_29);
R1IN_ADD_1_0_AXB_28_Z7492: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(28),
  I1 => R1IN_3(28),
  LO => R1IN_ADD_1_0_AXB_28);
R1IN_ADD_1_0_AXB_27_Z7493: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(27),
  I1 => R1IN_3(27),
  LO => R1IN_ADD_1_0_AXB_27);
R1IN_ADD_1_0_AXB_26_Z7494: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(26),
  I1 => R1IN_3(26),
  LO => R1IN_ADD_1_0_AXB_26);
R1IN_ADD_1_0_AXB_25_Z7495: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(25),
  I1 => R1IN_3(25),
  LO => R1IN_ADD_1_0_AXB_25);
R1IN_ADD_1_0_AXB_24_Z7496: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(24),
  I1 => R1IN_3(24),
  LO => R1IN_ADD_1_0_AXB_24);
R1IN_ADD_1_0_AXB_23_Z7497: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(23),
  I1 => R1IN_3(23),
  LO => R1IN_ADD_1_0_AXB_23);
R1IN_ADD_1_0_AXB_22_Z7498: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(22),
  I1 => R1IN_3(22),
  LO => R1IN_ADD_1_0_AXB_22);
R1IN_ADD_1_0_AXB_21_Z7499: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(21),
  I1 => R1IN_3(21),
  LO => R1IN_ADD_1_0_AXB_21);
R1IN_ADD_1_0_AXB_20_Z7500: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(20),
  I1 => R1IN_3(20),
  LO => R1IN_ADD_1_0_AXB_20);
R1IN_ADD_1_0_AXB_19_Z7501: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(19),
  I1 => R1IN_3(19),
  LO => R1IN_ADD_1_0_AXB_19);
R1IN_ADD_1_0_AXB_18_Z7502: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2(18),
  I1 => R1IN_3(18),
  LO => R1IN_ADD_1_0_AXB_18);
R1IN_ADD_1_0_AXB_16_Z7503: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F(16),
  I1 => R1IN_3F(16),
  LO => R1IN_ADD_1_0_AXB_16);
R1IN_ADD_1_0_AXB_15_Z7504: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F(15),
  I1 => R1IN_3F(15),
  LO => R1IN_ADD_1_0_AXB_15);
R1IN_ADD_1_0_AXB_14_Z7505: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F(14),
  I1 => R1IN_3F(14),
  LO => R1IN_ADD_1_0_AXB_14);
R1IN_ADD_1_0_AXB_13_Z7506: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F(13),
  I1 => R1IN_3F(13),
  LO => R1IN_ADD_1_0_AXB_13);
R1IN_ADD_1_0_AXB_12_Z7507: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F(12),
  I1 => R1IN_3F(12),
  LO => R1IN_ADD_1_0_AXB_12);
R1IN_ADD_1_0_AXB_11_Z7508: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F(11),
  I1 => R1IN_3F(11),
  LO => R1IN_ADD_1_0_AXB_11);
R1IN_ADD_1_0_AXB_10_Z7509: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F(10),
  I1 => R1IN_3F(10),
  LO => R1IN_ADD_1_0_AXB_10);
R1IN_ADD_1_0_AXB_9_Z7510: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F(9),
  I1 => R1IN_3F(9),
  LO => R1IN_ADD_1_0_AXB_9);
R1IN_ADD_1_0_AXB_8_Z7511: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F(8),
  I1 => R1IN_3F(8),
  LO => R1IN_ADD_1_0_AXB_8);
R1IN_ADD_1_0_AXB_7_Z7512: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F(7),
  I1 => R1IN_3F(7),
  LO => R1IN_ADD_1_0_AXB_7);
R1IN_ADD_1_0_AXB_6_Z7513: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F(6),
  I1 => R1IN_3F(6),
  LO => R1IN_ADD_1_0_AXB_6);
R1IN_ADD_1_0_AXB_5_Z7514: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F(5),
  I1 => R1IN_3F(5),
  LO => R1IN_ADD_1_0_AXB_5);
R1IN_ADD_1_0_AXB_4_Z7515: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F(4),
  I1 => R1IN_3F(4),
  LO => R1IN_ADD_1_0_AXB_4);
R1IN_ADD_1_0_AXB_3_Z7516: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F(3),
  I1 => R1IN_3F(3),
  LO => R1IN_ADD_1_0_AXB_3);
R1IN_ADD_1_0_AXB_2_Z7517: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F(2),
  I1 => R1IN_3F(2),
  LO => R1IN_ADD_1_0_AXB_2);
R1IN_ADD_1_0_AXB_1_Z7518: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F(1),
  I1 => R1IN_3F(1),
  LO => R1IN_ADD_1_0_AXB_1);
R1IN_ADD_1_0_AXB_0: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_2F(0),
  I1 => R1IN_3F(0),
  O => R1IN_ADD_1(0));
R1IN_ADD_2_0_AXB_0: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_ADD_1FF(0),
  I1 => R1IN_ADD_2_0,
  O => NN_11);
R1IN_4_ADD_2_1_AXB_34_Z7521: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(53),
  LO => R1IN_4_ADD_2_1_AXB_34);
R1IN_4_ADD_2_1_AXB_33_Z7522: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(52),
  LO => R1IN_4_ADD_2_1_AXB_33);
R1IN_4_ADD_2_1_AXB_32_Z7523: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(51),
  LO => R1IN_4_ADD_2_1_AXB_32);
R1IN_4_ADD_2_1_AXB_31_Z7524: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(50),
  LO => R1IN_4_ADD_2_1_AXB_31);
R1IN_4_ADD_2_1_AXB_30_Z7525: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(49),
  LO => R1IN_4_ADD_2_1_AXB_30);
R1IN_4_ADD_2_1_AXB_29_Z7526: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(48),
  LO => R1IN_4_ADD_2_1_AXB_29);
R1IN_4_ADD_2_1_AXB_28_Z7527: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(47),
  LO => R1IN_4_ADD_2_1_AXB_28);
R1IN_4_ADD_2_1_AXB_27_Z7528: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(46),
  LO => R1IN_4_ADD_2_1_AXB_27);
R1IN_4_ADD_2_1_AXB_26_Z7529: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(45),
  LO => R1IN_4_ADD_2_1_AXB_26);
R1IN_4_ADD_2_1_AXB_25_Z7530: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(44),
  LO => R1IN_4_ADD_2_1_AXB_25);
R1IN_4_ADD_2_1_AXB_24_Z7531: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(43),
  LO => R1IN_4_ADD_2_1_AXB_24);
R1IN_4_ADD_2_1_AXB_23_Z7532: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(42),
  LO => R1IN_4_ADD_2_1_AXB_23);
R1IN_4_ADD_2_1_AXB_22_Z7533: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(41),
  LO => R1IN_4_ADD_2_1_AXB_22);
R1IN_4_ADD_2_1_AXB_21_Z7534: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(40),
  LO => R1IN_4_ADD_2_1_AXB_21);
R1IN_4_ADD_2_1_AXB_20_Z7535: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(39),
  LO => R1IN_4_ADD_2_1_AXB_20);
R1IN_4_ADD_2_1_AXB_19_Z7536: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(38),
  LO => R1IN_4_ADD_2_1_AXB_19);
R1IN_4_ADD_2_1_AXB_18_Z7537: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(37),
  LO => R1IN_4_ADD_2_1_AXB_18);
R1IN_4_ADD_2_1_AXB_17_Z7538: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(36),
  LO => R1IN_4_ADD_2_1_AXB_17);
R1IN_4_ADD_2_1_AXB_16_Z7539: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(35),
  LO => R1IN_4_ADD_2_1_AXB_16);
R1IN_4_ADD_2_1_AXB_15_Z7540: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(34),
  LO => R1IN_4_ADD_2_1_AXB_15);
R1IN_4_ADD_2_1_AXB_14_Z7541: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(33),
  LO => R1IN_4_ADD_2_1_AXB_14);
R1IN_4_ADD_2_1_AXB_13_Z7542: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(32),
  LO => R1IN_4_ADD_2_1_AXB_13);
R1IN_4_ADD_2_1_AXB_12_Z7543: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(31),
  LO => R1IN_4_ADD_2_1_AXB_12);
R1IN_4_ADD_2_1_AXB_11_Z7544: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(30),
  LO => R1IN_4_ADD_2_1_AXB_11);
R1IN_4_ADD_2_1_AXB_10_Z7545: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(29),
  LO => R1IN_4_ADD_2_1_AXB_10);
R1IN_4_ADD_2_1_AXB_9_Z7546: LUT1_L 
generic map(
  INIT => X"2"
)
port map (
  I0 => R1IN_4_4(28),
  LO => R1IN_4_ADD_2_1_AXB_9);
R1IN_4_ADD_2_1_AXB_8_Z7547: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(27),
  I1 => NN_10,
  LO => R1IN_4_ADD_2_1_AXB_8);
R1IN_4_ADD_2_1_AXB_7_Z7548: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(26),
  I1 => NN_9,
  LO => R1IN_4_ADD_2_1_AXB_7);
R1IN_4_ADD_2_1_AXB_6_Z7549: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(25),
  I1 => NN_8,
  LO => R1IN_4_ADD_2_1_AXB_6);
R1IN_4_ADD_2_1_AXB_5_Z7550: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(24),
  I1 => NN_7,
  LO => R1IN_4_ADD_2_1_AXB_5);
R1IN_4_ADD_2_1_AXB_4_Z7551: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(23),
  I1 => NN_6,
  LO => R1IN_4_ADD_2_1_AXB_4);
R1IN_4_ADD_2_1_AXB_3_Z7552: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(22),
  I1 => NN_5,
  LO => R1IN_4_ADD_2_1_AXB_3);
R1IN_4_ADD_2_1_AXB_2_Z7553: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(21),
  I1 => NN_4,
  LO => R1IN_4_ADD_2_1_AXB_2);
R1IN_4_ADD_2_1_AXB_1_Z7554: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(20),
  I1 => NN_3,
  LO => R1IN_4_ADD_2_1_AXB_1);
R1IN_4_ADD_2_1_AXB_0_Z7555: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(19),
  I1 => R1IN_4_ADD_2_1,
  O => R1IN_4_ADD_2_1_AXB_0_RETI);
R1IN_4_ADD_2_0_AXB_35_Z7556: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4(18),
  I1 => R1IN_4_ADD_1(35),
  LO => R1IN_4_ADD_2_0_AXB_35);
R1IN_4_ADD_2_0_AXB_33_Z7557: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F(16),
  I1 => R1IN_4_ADD_1(33),
  LO => R1IN_4_ADD_2_0_AXB_33);
R1IN_4_ADD_2_0_AXB_32_Z7558: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F(15),
  I1 => R1IN_4_ADD_1(32),
  LO => R1IN_4_ADD_2_0_AXB_32);
R1IN_4_ADD_2_0_AXB_31_Z7559: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F(14),
  I1 => R1IN_4_ADD_1(31),
  LO => R1IN_4_ADD_2_0_AXB_31);
R1IN_4_ADD_2_0_AXB_30_Z7560: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F(13),
  I1 => R1IN_4_ADD_1(30),
  LO => R1IN_4_ADD_2_0_AXB_30);
R1IN_4_ADD_2_0_AXB_29_Z7561: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F(12),
  I1 => R1IN_4_ADD_1(29),
  LO => R1IN_4_ADD_2_0_AXB_29);
R1IN_4_ADD_2_0_AXB_28_Z7562: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F(11),
  I1 => R1IN_4_ADD_1(28),
  LO => R1IN_4_ADD_2_0_AXB_28);
R1IN_4_ADD_2_0_AXB_27_Z7563: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F(10),
  I1 => R1IN_4_ADD_1(27),
  LO => R1IN_4_ADD_2_0_AXB_27);
R1IN_4_ADD_2_0_AXB_26_Z7564: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F(9),
  I1 => R1IN_4_ADD_1(26),
  LO => R1IN_4_ADD_2_0_AXB_26);
R1IN_4_ADD_2_0_AXB_25_Z7565: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F(8),
  I1 => R1IN_4_ADD_1(25),
  LO => R1IN_4_ADD_2_0_AXB_25);
R1IN_4_ADD_2_0_AXB_24_Z7566: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F(7),
  I1 => R1IN_4_ADD_1(24),
  LO => R1IN_4_ADD_2_0_AXB_24);
R1IN_4_ADD_2_0_AXB_23_Z7567: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F(6),
  I1 => R1IN_4_ADD_1(23),
  LO => R1IN_4_ADD_2_0_AXB_23);
R1IN_4_ADD_2_0_AXB_22_Z7568: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F(5),
  I1 => R1IN_4_ADD_1(22),
  LO => R1IN_4_ADD_2_0_AXB_22);
R1IN_4_ADD_2_0_AXB_21_Z7569: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F(4),
  I1 => R1IN_4_ADD_1(21),
  LO => R1IN_4_ADD_2_0_AXB_21);
R1IN_4_ADD_2_0_AXB_20_Z7570: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F(3),
  I1 => R1IN_4_ADD_1(20),
  LO => R1IN_4_ADD_2_0_AXB_20);
R1IN_4_ADD_2_0_AXB_19_Z7571: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F(2),
  I1 => R1IN_4_ADD_1(19),
  LO => R1IN_4_ADD_2_0_AXB_19);
R1IN_4_ADD_2_0_AXB_18_Z7572: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F(1),
  I1 => R1IN_4_ADD_1(18),
  LO => R1IN_4_ADD_2_0_AXB_18);
R1IN_4_ADD_2_0_AXB_17_Z7573: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_4F(0),
  I1 => R1IN_4_ADD_1(17),
  LO => R1IN_4_ADD_2_0_AXB_17);
R1IN_4_ADD_2_0_AXB_16_Z7574: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F(33),
  I1 => R1IN_4_ADD_1(16),
  LO => R1IN_4_ADD_2_0_AXB_16);
R1IN_4_ADD_2_0_AXB_15_Z7575: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F(32),
  I1 => R1IN_4_ADD_1(15),
  LO => R1IN_4_ADD_2_0_AXB_15);
R1IN_4_ADD_2_0_AXB_14_Z7576: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F(31),
  I1 => R1IN_4_ADD_1(14),
  LO => R1IN_4_ADD_2_0_AXB_14);
R1IN_4_ADD_2_0_AXB_13_Z7577: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F(30),
  I1 => R1IN_4_ADD_1(13),
  LO => R1IN_4_ADD_2_0_AXB_13);
R1IN_4_ADD_2_0_AXB_12_Z7578: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F(29),
  I1 => R1IN_4_ADD_1(12),
  LO => R1IN_4_ADD_2_0_AXB_12);
R1IN_4_ADD_2_0_AXB_11_Z7579: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F(28),
  I1 => R1IN_4_ADD_1(11),
  LO => R1IN_4_ADD_2_0_AXB_11);
R1IN_4_ADD_2_0_AXB_10_Z7580: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F(27),
  I1 => R1IN_4_ADD_1(10),
  LO => R1IN_4_ADD_2_0_AXB_10);
R1IN_4_ADD_2_0_AXB_9_Z7581: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F(26),
  I1 => R1IN_4_ADD_1(9),
  LO => R1IN_4_ADD_2_0_AXB_9);
R1IN_4_ADD_2_0_AXB_8_Z7582: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F(25),
  I1 => R1IN_4_ADD_1(8),
  LO => R1IN_4_ADD_2_0_AXB_8);
R1IN_4_ADD_2_0_AXB_7_Z7583: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F(24),
  I1 => R1IN_4_ADD_1(7),
  LO => R1IN_4_ADD_2_0_AXB_7);
R1IN_4_ADD_2_0_AXB_6_Z7584: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F(23),
  I1 => R1IN_4_ADD_1(6),
  LO => R1IN_4_ADD_2_0_AXB_6);
R1IN_4_ADD_2_0_AXB_5_Z7585: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F(22),
  I1 => R1IN_4_ADD_1(5),
  LO => R1IN_4_ADD_2_0_AXB_5);
R1IN_4_ADD_2_0_AXB_4_Z7586: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F(21),
  I1 => R1IN_4_ADD_1(4),
  LO => R1IN_4_ADD_2_0_AXB_4);
R1IN_4_ADD_2_0_AXB_3_Z7587: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F(20),
  I1 => R1IN_4_ADD_1(3),
  LO => R1IN_4_ADD_2_0_AXB_3);
R1IN_4_ADD_2_0_AXB_2_Z7588: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F(19),
  I1 => R1IN_4_ADD_1(2),
  LO => R1IN_4_ADD_2_0_AXB_2);
R1IN_4_ADD_2_0_AXB_1_Z7589: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F(18),
  I1 => R1IN_4_ADD_1(1),
  LO => R1IN_4_ADD_2_0_AXB_1);
R1IN_4_ADD_2_0_AXB_0: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => R1IN_4_1F(17),
  I1 => R1IN_4_ADD_2_0,
  O => R1IN_4(17));
R1IN_4_ADD_1_S_43: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_43,
    CI => R1IN_4_ADD_1_CRY_42,
    O => NN_9);
R1IN_4_ADD_1_CRY_43: MUXCY port map (
    DI => R1IN_4_2F(43),
    CI => R1IN_4_ADD_1_CRY_42,
    S => R1IN_4_ADD_1_AXB_43,
    O => NN_10);
R1IN_4_ADD_1_S_42: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_42,
    CI => R1IN_4_ADD_1_CRY_41,
    O => NN_8);
R1IN_4_ADD_1_CRY_42_Z7594: MUXCY_L port map (
    DI => R1IN_4_2F(42),
    CI => R1IN_4_ADD_1_CRY_41,
    S => R1IN_4_ADD_1_AXB_42,
    LO => R1IN_4_ADD_1_CRY_42);
R1IN_4_ADD_1_S_41: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_41,
    CI => R1IN_4_ADD_1_CRY_40,
    O => NN_7);
R1IN_4_ADD_1_CRY_41_Z7596: MUXCY_L port map (
    DI => R1IN_4_2F(41),
    CI => R1IN_4_ADD_1_CRY_40,
    S => R1IN_4_ADD_1_AXB_41,
    LO => R1IN_4_ADD_1_CRY_41);
R1IN_4_ADD_1_S_40: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_40,
    CI => R1IN_4_ADD_1_CRY_39,
    O => NN_6);
R1IN_4_ADD_1_CRY_40_Z7598: MUXCY_L port map (
    DI => R1IN_4_2F(40),
    CI => R1IN_4_ADD_1_CRY_39,
    S => R1IN_4_ADD_1_AXB_40,
    LO => R1IN_4_ADD_1_CRY_40);
R1IN_4_ADD_1_S_39: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_39,
    CI => R1IN_4_ADD_1_CRY_38,
    O => NN_5);
R1IN_4_ADD_1_CRY_39_Z7600: MUXCY_L port map (
    DI => R1IN_4_2F(39),
    CI => R1IN_4_ADD_1_CRY_38,
    S => R1IN_4_ADD_1_AXB_39,
    LO => R1IN_4_ADD_1_CRY_39);
R1IN_4_ADD_1_S_38: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_38,
    CI => R1IN_4_ADD_1_CRY_37,
    O => NN_4);
R1IN_4_ADD_1_CRY_38_Z7602: MUXCY_L port map (
    DI => R1IN_4_2F(38),
    CI => R1IN_4_ADD_1_CRY_37,
    S => R1IN_4_ADD_1_AXB_38,
    LO => R1IN_4_ADD_1_CRY_38);
R1IN_4_ADD_1_S_37: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_37,
    CI => R1IN_4_ADD_1_CRY_36,
    O => NN_3);
R1IN_4_ADD_1_CRY_37_Z7604: MUXCY_L port map (
    DI => R1IN_4_2F(37),
    CI => R1IN_4_ADD_1_CRY_36,
    S => R1IN_4_ADD_1_AXB_37,
    LO => R1IN_4_ADD_1_CRY_37);
R1IN_4_ADD_1_S_36: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_36,
    CI => R1IN_4_ADD_1_CRY_35,
    O => R1IN_4_ADD_2_1);
R1IN_4_ADD_1_CRY_36_Z7606: MUXCY_L port map (
    DI => R1IN_4_2F(36),
    CI => R1IN_4_ADD_1_CRY_35,
    S => R1IN_4_ADD_1_AXB_36,
    LO => R1IN_4_ADD_1_CRY_36);
R1IN_4_ADD_1_S_35: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_35,
    CI => R1IN_4_ADD_1_CRY_34,
    O => R1IN_4_ADD_1(35));
R1IN_4_ADD_1_CRY_35_Z7608: MUXCY_L port map (
    DI => R1IN_4_2F(35),
    CI => R1IN_4_ADD_1_CRY_34,
    S => R1IN_4_ADD_1_AXB_35,
    LO => R1IN_4_ADD_1_CRY_35);
R1IN_4_ADD_1_S_34: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_34,
    CI => R1IN_4_ADD_1_CRY_33,
    O => R1IN_4_ADD_1(34));
R1IN_4_ADD_1_CRY_34_Z7610: MUXCY_L port map (
    DI => R1IN_4_2F(34),
    CI => R1IN_4_ADD_1_CRY_33,
    S => R1IN_4_ADD_1_AXB_34,
    LO => R1IN_4_ADD_1_CRY_34);
R1IN_4_ADD_1_S_33: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_33,
    CI => R1IN_4_ADD_1_CRY_32,
    O => R1IN_4_ADD_1(33));
R1IN_4_ADD_1_CRY_33_Z7612: MUXCY_L port map (
    DI => R1IN_4_2F(33),
    CI => R1IN_4_ADD_1_CRY_32,
    S => R1IN_4_ADD_1_AXB_33,
    LO => R1IN_4_ADD_1_CRY_33);
R1IN_4_ADD_1_S_32: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_32,
    CI => R1IN_4_ADD_1_CRY_31,
    O => R1IN_4_ADD_1(32));
R1IN_4_ADD_1_CRY_32_Z7614: MUXCY_L port map (
    DI => R1IN_4_2F(32),
    CI => R1IN_4_ADD_1_CRY_31,
    S => R1IN_4_ADD_1_AXB_32,
    LO => R1IN_4_ADD_1_CRY_32);
R1IN_4_ADD_1_S_31: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_31,
    CI => R1IN_4_ADD_1_CRY_30,
    O => R1IN_4_ADD_1(31));
R1IN_4_ADD_1_CRY_31_Z7616: MUXCY_L port map (
    DI => R1IN_4_2F(31),
    CI => R1IN_4_ADD_1_CRY_30,
    S => R1IN_4_ADD_1_AXB_31,
    LO => R1IN_4_ADD_1_CRY_31);
R1IN_4_ADD_1_S_30: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_30,
    CI => R1IN_4_ADD_1_CRY_29,
    O => R1IN_4_ADD_1(30));
R1IN_4_ADD_1_CRY_30_Z7618: MUXCY_L port map (
    DI => R1IN_4_2F(30),
    CI => R1IN_4_ADD_1_CRY_29,
    S => R1IN_4_ADD_1_AXB_30,
    LO => R1IN_4_ADD_1_CRY_30);
R1IN_4_ADD_1_S_29: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_29,
    CI => R1IN_4_ADD_1_CRY_28,
    O => R1IN_4_ADD_1(29));
R1IN_4_ADD_1_CRY_29_Z7620: MUXCY_L port map (
    DI => R1IN_4_2F(29),
    CI => R1IN_4_ADD_1_CRY_28,
    S => R1IN_4_ADD_1_AXB_29,
    LO => R1IN_4_ADD_1_CRY_29);
R1IN_4_ADD_1_S_28: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_28,
    CI => R1IN_4_ADD_1_CRY_27,
    O => R1IN_4_ADD_1(28));
R1IN_4_ADD_1_CRY_28_Z7622: MUXCY_L port map (
    DI => R1IN_4_2F(28),
    CI => R1IN_4_ADD_1_CRY_27,
    S => R1IN_4_ADD_1_AXB_28,
    LO => R1IN_4_ADD_1_CRY_28);
R1IN_4_ADD_1_S_27: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_27,
    CI => R1IN_4_ADD_1_CRY_26,
    O => R1IN_4_ADD_1(27));
R1IN_4_ADD_1_CRY_27_Z7624: MUXCY_L port map (
    DI => R1IN_4_2F(27),
    CI => R1IN_4_ADD_1_CRY_26,
    S => R1IN_4_ADD_1_AXB_27,
    LO => R1IN_4_ADD_1_CRY_27);
R1IN_4_ADD_1_S_26: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_26,
    CI => R1IN_4_ADD_1_CRY_25,
    O => R1IN_4_ADD_1(26));
R1IN_4_ADD_1_CRY_26_Z7626: MUXCY_L port map (
    DI => R1IN_4_2F(26),
    CI => R1IN_4_ADD_1_CRY_25,
    S => R1IN_4_ADD_1_AXB_26,
    LO => R1IN_4_ADD_1_CRY_26);
R1IN_4_ADD_1_S_25: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_25,
    CI => R1IN_4_ADD_1_CRY_24,
    O => R1IN_4_ADD_1(25));
R1IN_4_ADD_1_CRY_25_Z7628: MUXCY_L port map (
    DI => R1IN_4_2F(25),
    CI => R1IN_4_ADD_1_CRY_24,
    S => R1IN_4_ADD_1_AXB_25,
    LO => R1IN_4_ADD_1_CRY_25);
R1IN_4_ADD_1_S_24: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_24,
    CI => R1IN_4_ADD_1_CRY_23,
    O => R1IN_4_ADD_1(24));
R1IN_4_ADD_1_CRY_24_Z7630: MUXCY_L port map (
    DI => R1IN_4_2F(24),
    CI => R1IN_4_ADD_1_CRY_23,
    S => R1IN_4_ADD_1_AXB_24,
    LO => R1IN_4_ADD_1_CRY_24);
R1IN_4_ADD_1_S_23: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_23,
    CI => R1IN_4_ADD_1_CRY_22,
    O => R1IN_4_ADD_1(23));
R1IN_4_ADD_1_CRY_23_Z7632: MUXCY_L port map (
    DI => R1IN_4_2F(23),
    CI => R1IN_4_ADD_1_CRY_22,
    S => R1IN_4_ADD_1_AXB_23,
    LO => R1IN_4_ADD_1_CRY_23);
R1IN_4_ADD_1_S_22: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_22,
    CI => R1IN_4_ADD_1_CRY_21,
    O => R1IN_4_ADD_1(22));
R1IN_4_ADD_1_CRY_22_Z7634: MUXCY_L port map (
    DI => R1IN_4_2F(22),
    CI => R1IN_4_ADD_1_CRY_21,
    S => R1IN_4_ADD_1_AXB_22,
    LO => R1IN_4_ADD_1_CRY_22);
R1IN_4_ADD_1_S_21: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_21,
    CI => R1IN_4_ADD_1_CRY_20,
    O => R1IN_4_ADD_1(21));
R1IN_4_ADD_1_CRY_21_Z7636: MUXCY_L port map (
    DI => R1IN_4_2F(21),
    CI => R1IN_4_ADD_1_CRY_20,
    S => R1IN_4_ADD_1_AXB_21,
    LO => R1IN_4_ADD_1_CRY_21);
R1IN_4_ADD_1_S_20: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_20,
    CI => R1IN_4_ADD_1_CRY_19,
    O => R1IN_4_ADD_1(20));
R1IN_4_ADD_1_CRY_20_Z7638: MUXCY_L port map (
    DI => R1IN_4_2F(20),
    CI => R1IN_4_ADD_1_CRY_19,
    S => R1IN_4_ADD_1_AXB_20,
    LO => R1IN_4_ADD_1_CRY_20);
R1IN_4_ADD_1_S_19: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_19,
    CI => R1IN_4_ADD_1_CRY_18,
    O => R1IN_4_ADD_1(19));
R1IN_4_ADD_1_CRY_19_Z7640: MUXCY_L port map (
    DI => R1IN_4_2F(19),
    CI => R1IN_4_ADD_1_CRY_18,
    S => R1IN_4_ADD_1_AXB_19,
    LO => R1IN_4_ADD_1_CRY_19);
R1IN_4_ADD_1_S_18: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_18,
    CI => R1IN_4_ADD_1_CRY_17,
    O => R1IN_4_ADD_1(18));
R1IN_4_ADD_1_CRY_18_Z7642: MUXCY_L port map (
    DI => R1IN_4_2F(18),
    CI => R1IN_4_ADD_1_CRY_17,
    S => R1IN_4_ADD_1_AXB_18,
    LO => R1IN_4_ADD_1_CRY_18);
R1IN_4_ADD_1_S_17: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_17,
    CI => R1IN_4_ADD_1_CRY_16,
    O => R1IN_4_ADD_1(17));
R1IN_4_ADD_1_CRY_17_Z7644: MUXCY_L port map (
    DI => R1IN_4_2F(17),
    CI => R1IN_4_ADD_1_CRY_16,
    S => R1IN_4_ADD_1_AXB_17,
    LO => R1IN_4_ADD_1_CRY_17);
R1IN_4_ADD_1_S_16: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_16,
    CI => R1IN_4_ADD_1_CRY_15,
    O => R1IN_4_ADD_1(16));
R1IN_4_ADD_1_CRY_16_Z7646: MUXCY_L port map (
    DI => R1IN_4_2F(16),
    CI => R1IN_4_ADD_1_CRY_15,
    S => R1IN_4_ADD_1_AXB_16,
    LO => R1IN_4_ADD_1_CRY_16);
R1IN_4_ADD_1_S_15: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_15,
    CI => R1IN_4_ADD_1_CRY_14,
    O => R1IN_4_ADD_1(15));
R1IN_4_ADD_1_CRY_15_Z7648: MUXCY_L port map (
    DI => R1IN_4_2F(15),
    CI => R1IN_4_ADD_1_CRY_14,
    S => R1IN_4_ADD_1_AXB_15,
    LO => R1IN_4_ADD_1_CRY_15);
R1IN_4_ADD_1_S_14: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_14,
    CI => R1IN_4_ADD_1_CRY_13,
    O => R1IN_4_ADD_1(14));
R1IN_4_ADD_1_CRY_14_Z7650: MUXCY_L port map (
    DI => R1IN_4_2F(14),
    CI => R1IN_4_ADD_1_CRY_13,
    S => R1IN_4_ADD_1_AXB_14,
    LO => R1IN_4_ADD_1_CRY_14);
R1IN_4_ADD_1_S_13: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_13,
    CI => R1IN_4_ADD_1_CRY_12,
    O => R1IN_4_ADD_1(13));
R1IN_4_ADD_1_CRY_13_Z7652: MUXCY_L port map (
    DI => R1IN_4_2F(13),
    CI => R1IN_4_ADD_1_CRY_12,
    S => R1IN_4_ADD_1_AXB_13,
    LO => R1IN_4_ADD_1_CRY_13);
R1IN_4_ADD_1_S_12: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_12,
    CI => R1IN_4_ADD_1_CRY_11,
    O => R1IN_4_ADD_1(12));
R1IN_4_ADD_1_CRY_12_Z7654: MUXCY_L port map (
    DI => R1IN_4_2F(12),
    CI => R1IN_4_ADD_1_CRY_11,
    S => R1IN_4_ADD_1_AXB_12,
    LO => R1IN_4_ADD_1_CRY_12);
R1IN_4_ADD_1_S_11: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_11,
    CI => R1IN_4_ADD_1_CRY_10,
    O => R1IN_4_ADD_1(11));
R1IN_4_ADD_1_CRY_11_Z7656: MUXCY_L port map (
    DI => R1IN_4_2F(11),
    CI => R1IN_4_ADD_1_CRY_10,
    S => R1IN_4_ADD_1_AXB_11,
    LO => R1IN_4_ADD_1_CRY_11);
R1IN_4_ADD_1_S_10: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_10,
    CI => R1IN_4_ADD_1_CRY_9,
    O => R1IN_4_ADD_1(10));
R1IN_4_ADD_1_CRY_10_Z7658: MUXCY_L port map (
    DI => R1IN_4_2F(10),
    CI => R1IN_4_ADD_1_CRY_9,
    S => R1IN_4_ADD_1_AXB_10,
    LO => R1IN_4_ADD_1_CRY_10);
R1IN_4_ADD_1_S_9: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_9,
    CI => R1IN_4_ADD_1_CRY_8,
    O => R1IN_4_ADD_1(9));
R1IN_4_ADD_1_CRY_9_Z7660: MUXCY_L port map (
    DI => R1IN_4_2F(9),
    CI => R1IN_4_ADD_1_CRY_8,
    S => R1IN_4_ADD_1_AXB_9,
    LO => R1IN_4_ADD_1_CRY_9);
R1IN_4_ADD_1_S_8: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_8,
    CI => R1IN_4_ADD_1_CRY_7,
    O => R1IN_4_ADD_1(8));
R1IN_4_ADD_1_CRY_8_Z7662: MUXCY_L port map (
    DI => R1IN_4_2F(8),
    CI => R1IN_4_ADD_1_CRY_7,
    S => R1IN_4_ADD_1_AXB_8,
    LO => R1IN_4_ADD_1_CRY_8);
R1IN_4_ADD_1_S_7: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_7,
    CI => R1IN_4_ADD_1_CRY_6,
    O => R1IN_4_ADD_1(7));
R1IN_4_ADD_1_CRY_7_Z7664: MUXCY_L port map (
    DI => R1IN_4_2F(7),
    CI => R1IN_4_ADD_1_CRY_6,
    S => R1IN_4_ADD_1_AXB_7,
    LO => R1IN_4_ADD_1_CRY_7);
R1IN_4_ADD_1_S_6: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_6,
    CI => R1IN_4_ADD_1_CRY_5,
    O => R1IN_4_ADD_1(6));
R1IN_4_ADD_1_CRY_6_Z7666: MUXCY_L port map (
    DI => R1IN_4_2F(6),
    CI => R1IN_4_ADD_1_CRY_5,
    S => R1IN_4_ADD_1_AXB_6,
    LO => R1IN_4_ADD_1_CRY_6);
R1IN_4_ADD_1_S_5: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_5,
    CI => R1IN_4_ADD_1_CRY_4,
    O => R1IN_4_ADD_1(5));
R1IN_4_ADD_1_CRY_5_Z7668: MUXCY_L port map (
    DI => R1IN_4_2F(5),
    CI => R1IN_4_ADD_1_CRY_4,
    S => R1IN_4_ADD_1_AXB_5,
    LO => R1IN_4_ADD_1_CRY_5);
R1IN_4_ADD_1_S_4: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_4,
    CI => R1IN_4_ADD_1_CRY_3,
    O => R1IN_4_ADD_1(4));
R1IN_4_ADD_1_CRY_4_Z7670: MUXCY_L port map (
    DI => R1IN_4_2F(4),
    CI => R1IN_4_ADD_1_CRY_3,
    S => R1IN_4_ADD_1_AXB_4,
    LO => R1IN_4_ADD_1_CRY_4);
R1IN_4_ADD_1_S_3: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_3,
    CI => R1IN_4_ADD_1_CRY_2,
    O => R1IN_4_ADD_1(3));
R1IN_4_ADD_1_CRY_3_Z7672: MUXCY_L port map (
    DI => R1IN_4_2F(3),
    CI => R1IN_4_ADD_1_CRY_2,
    S => R1IN_4_ADD_1_AXB_3,
    LO => R1IN_4_ADD_1_CRY_3);
R1IN_4_ADD_1_S_2: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_2,
    CI => R1IN_4_ADD_1_CRY_1,
    O => R1IN_4_ADD_1(2));
R1IN_4_ADD_1_CRY_2_Z7674: MUXCY_L port map (
    DI => R1IN_4_2F(2),
    CI => R1IN_4_ADD_1_CRY_1,
    S => R1IN_4_ADD_1_AXB_2,
    LO => R1IN_4_ADD_1_CRY_2);
R1IN_4_ADD_1_S_1: XORCY port map (
    LI => R1IN_4_ADD_1_AXB_1,
    CI => R1IN_4_ADD_1_CRY_0,
    O => R1IN_4_ADD_1(1));
R1IN_4_ADD_1_CRY_1_Z7676: MUXCY_L port map (
    DI => R1IN_4_2F(1),
    CI => R1IN_4_ADD_1_CRY_0,
    S => R1IN_4_ADD_1_AXB_1,
    LO => R1IN_4_ADD_1_CRY_1);
R1IN_4_ADD_1_CRY_0_Z7677: MUXCY_L port map (
    DI => NN_12,
    CI => NN_1,
    S => R1IN_4_ADD_2_0,
    LO => R1IN_4_ADD_1_CRY_0);
R1IN_4_4_ADD_2_S_36: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_36,
    CI => R1IN_4_4_ADD_2_CRY_35,
    O => R1IN_4_4(53));
R1IN_4_4_ADD_2_S_35: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_35,
    CI => R1IN_4_4_ADD_2_CRY_34,
    O => R1IN_4_4(52));
R1IN_4_4_ADD_2_CRY_35_Z7680: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_4_ADD_2_CRY_34,
    S => R1IN_4_4_ADD_2_AXB_35,
    LO => R1IN_4_4_ADD_2_CRY_35);
R1IN_4_4_ADD_2_S_34: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_34,
    CI => R1IN_4_4_ADD_2_CRY_33,
    O => R1IN_4_4(51));
R1IN_4_4_ADD_2_CRY_34_Z7682: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_4_ADD_2_CRY_33,
    S => R1IN_4_4_ADD_2_AXB_34,
    LO => R1IN_4_4_ADD_2_CRY_34);
R1IN_4_4_ADD_2_S_33: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_33,
    CI => R1IN_4_4_ADD_2_CRY_32,
    O => R1IN_4_4(50));
R1IN_4_4_ADD_2_CRY_33_Z7684: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_4_ADD_2_CRY_32,
    S => R1IN_4_4_ADD_2_AXB_33,
    LO => R1IN_4_4_ADD_2_CRY_33);
R1IN_4_4_ADD_2_S_32: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_32,
    CI => R1IN_4_4_ADD_2_CRY_31,
    O => R1IN_4_4(49));
R1IN_4_4_ADD_2_CRY_32_Z7686: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_4_ADD_2_CRY_31,
    S => R1IN_4_4_ADD_2_AXB_32,
    LO => R1IN_4_4_ADD_2_CRY_32);
R1IN_4_4_ADD_2_S_31: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_31,
    CI => R1IN_4_4_ADD_2_CRY_30,
    O => R1IN_4_4(48));
R1IN_4_4_ADD_2_CRY_31_Z7688: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_4_ADD_2_CRY_30,
    S => R1IN_4_4_ADD_2_AXB_31,
    LO => R1IN_4_4_ADD_2_CRY_31);
R1IN_4_4_ADD_2_S_30: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_30,
    CI => R1IN_4_4_ADD_2_CRY_29,
    O => R1IN_4_4(47));
R1IN_4_4_ADD_2_CRY_30_Z7690: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_4_ADD_2_CRY_29,
    S => R1IN_4_4_ADD_2_AXB_30,
    LO => R1IN_4_4_ADD_2_CRY_30);
R1IN_4_4_ADD_2_S_29: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_29,
    CI => R1IN_4_4_ADD_2_CRY_28,
    O => R1IN_4_4(46));
R1IN_4_4_ADD_2_CRY_29_Z7692: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_4_ADD_2_CRY_28,
    S => R1IN_4_4_ADD_2_AXB_29,
    LO => R1IN_4_4_ADD_2_CRY_29);
R1IN_4_4_ADD_2_S_28: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_28,
    CI => R1IN_4_4_ADD_2_CRY_27,
    O => R1IN_4_4(45));
R1IN_4_4_ADD_2_CRY_28_Z7694: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_4_ADD_2_CRY_27,
    S => R1IN_4_4_ADD_2_AXB_28,
    LO => R1IN_4_4_ADD_2_CRY_28);
R1IN_4_4_ADD_2_S_27: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_27,
    CI => R1IN_4_4_ADD_2_CRY_26,
    O => R1IN_4_4(44));
R1IN_4_4_ADD_2_CRY_27_Z7696: MUXCY_L port map (
    DI => R1IN_4_4_4F(10),
    CI => R1IN_4_4_ADD_2_CRY_26,
    S => R1IN_4_4_ADD_2_AXB_27,
    LO => R1IN_4_4_ADD_2_CRY_27);
R1IN_4_4_ADD_2_S_26: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_26,
    CI => R1IN_4_4_ADD_2_CRY_25,
    O => R1IN_4_4(43));
R1IN_4_4_ADD_2_CRY_26_Z7698: MUXCY_L port map (
    DI => R1IN_4_4_4F(9),
    CI => R1IN_4_4_ADD_2_CRY_25,
    S => R1IN_4_4_ADD_2_AXB_26,
    LO => R1IN_4_4_ADD_2_CRY_26);
R1IN_4_4_ADD_2_S_25: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_25,
    CI => R1IN_4_4_ADD_2_CRY_24,
    O => R1IN_4_4(42));
R1IN_4_4_ADD_2_CRY_25_Z7700: MUXCY_L port map (
    DI => R1IN_4_4_4F(8),
    CI => R1IN_4_4_ADD_2_CRY_24,
    S => R1IN_4_4_ADD_2_AXB_25,
    LO => R1IN_4_4_ADD_2_CRY_25);
R1IN_4_4_ADD_2_S_24: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_24,
    CI => R1IN_4_4_ADD_2_CRY_23,
    O => R1IN_4_4(41));
R1IN_4_4_ADD_2_CRY_24_Z7702: MUXCY_L port map (
    DI => R1IN_4_4_4F(7),
    CI => R1IN_4_4_ADD_2_CRY_23,
    S => R1IN_4_4_ADD_2_AXB_24,
    LO => R1IN_4_4_ADD_2_CRY_24);
R1IN_4_4_ADD_2_S_23: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_23,
    CI => R1IN_4_4_ADD_2_CRY_22,
    O => R1IN_4_4(40));
R1IN_4_4_ADD_2_CRY_23_Z7704: MUXCY_L port map (
    DI => R1IN_4_4_4F(6),
    CI => R1IN_4_4_ADD_2_CRY_22,
    S => R1IN_4_4_ADD_2_AXB_23,
    LO => R1IN_4_4_ADD_2_CRY_23);
R1IN_4_4_ADD_2_S_22: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_22,
    CI => R1IN_4_4_ADD_2_CRY_21,
    O => R1IN_4_4(39));
R1IN_4_4_ADD_2_CRY_22_Z7706: MUXCY_L port map (
    DI => R1IN_4_4_4F(5),
    CI => R1IN_4_4_ADD_2_CRY_21,
    S => R1IN_4_4_ADD_2_AXB_22,
    LO => R1IN_4_4_ADD_2_CRY_22);
R1IN_4_4_ADD_2_S_21: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_21,
    CI => R1IN_4_4_ADD_2_CRY_20,
    O => R1IN_4_4(38));
R1IN_4_4_ADD_2_CRY_21_Z7708: MUXCY_L port map (
    DI => R1IN_4_4_4F(4),
    CI => R1IN_4_4_ADD_2_CRY_20,
    S => R1IN_4_4_ADD_2_AXB_21,
    LO => R1IN_4_4_ADD_2_CRY_21);
R1IN_4_4_ADD_2_S_20: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_20,
    CI => R1IN_4_4_ADD_2_CRY_19,
    O => R1IN_4_4(37));
R1IN_4_4_ADD_2_CRY_20_Z7710: MUXCY_L port map (
    DI => R1IN_4_4_4F(3),
    CI => R1IN_4_4_ADD_2_CRY_19,
    S => R1IN_4_4_ADD_2_AXB_20,
    LO => R1IN_4_4_ADD_2_CRY_20);
R1IN_4_4_ADD_2_S_19: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_19,
    CI => R1IN_4_4_ADD_2_CRY_18,
    O => R1IN_4_4(36));
R1IN_4_4_ADD_2_CRY_19_Z7712: MUXCY_L port map (
    DI => R1IN_4_4_4F(2),
    CI => R1IN_4_4_ADD_2_CRY_18,
    S => R1IN_4_4_ADD_2_AXB_19,
    LO => R1IN_4_4_ADD_2_CRY_19);
R1IN_4_4_ADD_2_S_18: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_18,
    CI => R1IN_4_4_ADD_2_CRY_17,
    O => R1IN_4_4(35));
R1IN_4_4_ADD_2_CRY_18_Z7714: MUXCY_L port map (
    DI => R1IN_4_4_4F(1),
    CI => R1IN_4_4_ADD_2_CRY_17,
    S => R1IN_4_4_ADD_2_AXB_18,
    LO => R1IN_4_4_ADD_2_CRY_18);
R1IN_4_4_ADD_2_S_17: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_17,
    CI => R1IN_4_4_ADD_2_CRY_16,
    O => R1IN_4_4(34));
R1IN_4_4_ADD_2_CRY_17_Z7716: MUXCY_L port map (
    DI => R1IN_4_4_4F(0),
    CI => R1IN_4_4_ADD_2_CRY_16,
    S => R1IN_4_4_ADD_2_AXB_17,
    LO => R1IN_4_4_ADD_2_CRY_17);
R1IN_4_4_ADD_2_S_16: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_16,
    CI => R1IN_4_4_ADD_2_CRY_15,
    O => R1IN_4_4(33));
R1IN_4_4_ADD_2_CRY_16_Z7718: MUXCY_L port map (
    DI => R1IN_4_4_1F(33),
    CI => R1IN_4_4_ADD_2_CRY_15,
    S => R1IN_4_4_ADD_2_AXB_16,
    LO => R1IN_4_4_ADD_2_CRY_16);
R1IN_4_4_ADD_2_S_15: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_15,
    CI => R1IN_4_4_ADD_2_CRY_14,
    O => R1IN_4_4(32));
R1IN_4_4_ADD_2_CRY_15_Z7720: MUXCY_L port map (
    DI => R1IN_4_4_1F(32),
    CI => R1IN_4_4_ADD_2_CRY_14,
    S => R1IN_4_4_ADD_2_AXB_15,
    LO => R1IN_4_4_ADD_2_CRY_15);
R1IN_4_4_ADD_2_S_14: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_14,
    CI => R1IN_4_4_ADD_2_CRY_13,
    O => R1IN_4_4(31));
R1IN_4_4_ADD_2_CRY_14_Z7722: MUXCY_L port map (
    DI => R1IN_4_4_1F(31),
    CI => R1IN_4_4_ADD_2_CRY_13,
    S => R1IN_4_4_ADD_2_AXB_14,
    LO => R1IN_4_4_ADD_2_CRY_14);
R1IN_4_4_ADD_2_S_13: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_13,
    CI => R1IN_4_4_ADD_2_CRY_12,
    O => R1IN_4_4(30));
R1IN_4_4_ADD_2_CRY_13_Z7724: MUXCY_L port map (
    DI => R1IN_4_4_1F(30),
    CI => R1IN_4_4_ADD_2_CRY_12,
    S => R1IN_4_4_ADD_2_AXB_13,
    LO => R1IN_4_4_ADD_2_CRY_13);
R1IN_4_4_ADD_2_S_12: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_12,
    CI => R1IN_4_4_ADD_2_CRY_11,
    O => R1IN_4_4(29));
R1IN_4_4_ADD_2_CRY_12_Z7726: MUXCY_L port map (
    DI => R1IN_4_4_1F(29),
    CI => R1IN_4_4_ADD_2_CRY_11,
    S => R1IN_4_4_ADD_2_AXB_12,
    LO => R1IN_4_4_ADD_2_CRY_12);
R1IN_4_4_ADD_2_S_11: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_11,
    CI => R1IN_4_4_ADD_2_CRY_10,
    O => R1IN_4_4(28));
R1IN_4_4_ADD_2_CRY_11_Z7728: MUXCY_L port map (
    DI => R1IN_4_4_1F(28),
    CI => R1IN_4_4_ADD_2_CRY_10,
    S => R1IN_4_4_ADD_2_AXB_11,
    LO => R1IN_4_4_ADD_2_CRY_11);
R1IN_4_4_ADD_2_S_10: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_10,
    CI => R1IN_4_4_ADD_2_CRY_9,
    O => R1IN_4_4(27));
R1IN_4_4_ADD_2_CRY_10_Z7730: MUXCY_L port map (
    DI => R1IN_4_4_1F(27),
    CI => R1IN_4_4_ADD_2_CRY_9,
    S => R1IN_4_4_ADD_2_AXB_10,
    LO => R1IN_4_4_ADD_2_CRY_10);
R1IN_4_4_ADD_2_S_9: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_9,
    CI => R1IN_4_4_ADD_2_CRY_8,
    O => R1IN_4_4(26));
R1IN_4_4_ADD_2_CRY_9_Z7732: MUXCY_L port map (
    DI => R1IN_4_4_1F(26),
    CI => R1IN_4_4_ADD_2_CRY_8,
    S => R1IN_4_4_ADD_2_AXB_9,
    LO => R1IN_4_4_ADD_2_CRY_9);
R1IN_4_4_ADD_2_S_8: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_8,
    CI => R1IN_4_4_ADD_2_CRY_7,
    O => R1IN_4_4(25));
R1IN_4_4_ADD_2_CRY_8_Z7734: MUXCY_L port map (
    DI => R1IN_4_4_1F(25),
    CI => R1IN_4_4_ADD_2_CRY_7,
    S => R1IN_4_4_ADD_2_AXB_8,
    LO => R1IN_4_4_ADD_2_CRY_8);
R1IN_4_4_ADD_2_S_7: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_7,
    CI => R1IN_4_4_ADD_2_CRY_6,
    O => R1IN_4_4(24));
R1IN_4_4_ADD_2_CRY_7_Z7736: MUXCY_L port map (
    DI => R1IN_4_4_1F(24),
    CI => R1IN_4_4_ADD_2_CRY_6,
    S => R1IN_4_4_ADD_2_AXB_7,
    LO => R1IN_4_4_ADD_2_CRY_7);
R1IN_4_4_ADD_2_S_6: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_6,
    CI => R1IN_4_4_ADD_2_CRY_5,
    O => R1IN_4_4(23));
R1IN_4_4_ADD_2_CRY_6_Z7738: MUXCY_L port map (
    DI => R1IN_4_4_1F(23),
    CI => R1IN_4_4_ADD_2_CRY_5,
    S => R1IN_4_4_ADD_2_AXB_6,
    LO => R1IN_4_4_ADD_2_CRY_6);
R1IN_4_4_ADD_2_S_5: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_5,
    CI => R1IN_4_4_ADD_2_CRY_4,
    O => R1IN_4_4(22));
R1IN_4_4_ADD_2_CRY_5_Z7740: MUXCY_L port map (
    DI => R1IN_4_4_1F(22),
    CI => R1IN_4_4_ADD_2_CRY_4,
    S => R1IN_4_4_ADD_2_AXB_5,
    LO => R1IN_4_4_ADD_2_CRY_5);
R1IN_4_4_ADD_2_S_4: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_4,
    CI => R1IN_4_4_ADD_2_CRY_3,
    O => R1IN_4_4(21));
R1IN_4_4_ADD_2_CRY_4_Z7742: MUXCY_L port map (
    DI => R1IN_4_4_1F(21),
    CI => R1IN_4_4_ADD_2_CRY_3,
    S => R1IN_4_4_ADD_2_AXB_4,
    LO => R1IN_4_4_ADD_2_CRY_4);
R1IN_4_4_ADD_2_S_3: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_3,
    CI => R1IN_4_4_ADD_2_CRY_2,
    O => R1IN_4_4(20));
R1IN_4_4_ADD_2_CRY_3_Z7744: MUXCY_L port map (
    DI => R1IN_4_4_1F(20),
    CI => R1IN_4_4_ADD_2_CRY_2,
    S => R1IN_4_4_ADD_2_AXB_3,
    LO => R1IN_4_4_ADD_2_CRY_3);
R1IN_4_4_ADD_2_S_2: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_2,
    CI => R1IN_4_4_ADD_2_CRY_1,
    O => R1IN_4_4(19));
R1IN_4_4_ADD_2_CRY_2_Z7746: MUXCY_L port map (
    DI => R1IN_4_4_1F(19),
    CI => R1IN_4_4_ADD_2_CRY_1,
    S => R1IN_4_4_ADD_2_AXB_2,
    LO => R1IN_4_4_ADD_2_CRY_2);
R1IN_4_4_ADD_2_S_1: XORCY port map (
    LI => R1IN_4_4_ADD_2_AXB_1,
    CI => R1IN_4_4_ADD_2_CRY_0,
    O => R1IN_4_4(18));
R1IN_4_4_ADD_2_CRY_1_Z7748: MUXCY_L port map (
    DI => R1IN_4_4_1F(18),
    CI => R1IN_4_4_ADD_2_CRY_0,
    S => R1IN_4_4_ADD_2_AXB_1,
    LO => R1IN_4_4_ADD_2_CRY_1);
R1IN_4_4_ADD_2_CRY_0_Z7749: MUXCY_L port map (
    DI => R1IN_4_4_ADD_2,
    CI => NN_1,
    S => R1IN_4_4(17),
    LO => R1IN_4_4_ADD_2_CRY_0);
R1IN_2_ADD_1_S_43: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_43,
    CI => R1IN_2_ADD_1_CRY_42,
    O => R1IN_2(60));
R1IN_2_ADD_1_S_42: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_42,
    CI => R1IN_2_ADD_1_CRY_41,
    O => R1IN_2(59));
R1IN_2_ADD_1_CRY_42_Z7752: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_41,
    S => R1IN_2_ADD_1_AXB_42,
    LO => R1IN_2_ADD_1_CRY_42);
R1IN_2_ADD_1_S_41: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_41,
    CI => R1IN_2_ADD_1_CRY_40,
    O => R1IN_2(58));
R1IN_2_ADD_1_CRY_41_Z7754: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_40,
    S => R1IN_2_ADD_1_AXB_41,
    LO => R1IN_2_ADD_1_CRY_41);
R1IN_2_ADD_1_S_40: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_40,
    CI => R1IN_2_ADD_1_CRY_39,
    O => R1IN_2(57));
R1IN_2_ADD_1_CRY_40_Z7756: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_39,
    S => R1IN_2_ADD_1_AXB_40,
    LO => R1IN_2_ADD_1_CRY_40);
R1IN_2_ADD_1_S_39: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_39,
    CI => R1IN_2_ADD_1_CRY_38,
    O => R1IN_2(56));
R1IN_2_ADD_1_CRY_39_Z7758: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_38,
    S => R1IN_2_ADD_1_AXB_39,
    LO => R1IN_2_ADD_1_CRY_39);
R1IN_2_ADD_1_S_38: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_38,
    CI => R1IN_2_ADD_1_CRY_37,
    O => R1IN_2(55));
R1IN_2_ADD_1_CRY_38_Z7760: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_37,
    S => R1IN_2_ADD_1_AXB_38,
    LO => R1IN_2_ADD_1_CRY_38);
R1IN_2_ADD_1_S_37: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_37,
    CI => R1IN_2_ADD_1_CRY_36,
    O => R1IN_2(54));
R1IN_2_ADD_1_CRY_37_Z7762: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_36,
    S => R1IN_2_ADD_1_AXB_37,
    LO => R1IN_2_ADD_1_CRY_37);
R1IN_2_ADD_1_S_36: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_36,
    CI => R1IN_2_ADD_1_CRY_35,
    O => R1IN_2(53));
R1IN_2_ADD_1_CRY_36_Z7764: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_35,
    S => R1IN_2_ADD_1_AXB_36,
    LO => R1IN_2_ADD_1_CRY_36);
R1IN_2_ADD_1_S_35: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_35,
    CI => R1IN_2_ADD_1_CRY_34,
    O => R1IN_2(52));
R1IN_2_ADD_1_CRY_35_Z7766: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_34,
    S => R1IN_2_ADD_1_AXB_35,
    LO => R1IN_2_ADD_1_CRY_35);
R1IN_2_ADD_1_S_34: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_34,
    CI => R1IN_2_ADD_1_CRY_33,
    O => R1IN_2(51));
R1IN_2_ADD_1_CRY_34_Z7768: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_33,
    S => R1IN_2_ADD_1_AXB_34,
    LO => R1IN_2_ADD_1_CRY_34);
R1IN_2_ADD_1_S_33: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_33,
    CI => R1IN_2_ADD_1_CRY_32,
    O => R1IN_2(50));
R1IN_2_ADD_1_CRY_33_Z7770: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_32,
    S => R1IN_2_ADD_1_AXB_33,
    LO => R1IN_2_ADD_1_CRY_33);
R1IN_2_ADD_1_S_32: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_32,
    CI => R1IN_2_ADD_1_CRY_31,
    O => R1IN_2(49));
R1IN_2_ADD_1_CRY_32_Z7772: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_31,
    S => R1IN_2_ADD_1_AXB_32,
    LO => R1IN_2_ADD_1_CRY_32);
R1IN_2_ADD_1_S_31: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_31,
    CI => R1IN_2_ADD_1_CRY_30,
    O => R1IN_2(48));
R1IN_2_ADD_1_CRY_31_Z7774: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_30,
    S => R1IN_2_ADD_1_AXB_31,
    LO => R1IN_2_ADD_1_CRY_31);
R1IN_2_ADD_1_S_30: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_30,
    CI => R1IN_2_ADD_1_CRY_29,
    O => R1IN_2(47));
R1IN_2_ADD_1_CRY_30_Z7776: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_29,
    S => R1IN_2_ADD_1_AXB_30,
    LO => R1IN_2_ADD_1_CRY_30);
R1IN_2_ADD_1_S_29: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_29,
    CI => R1IN_2_ADD_1_CRY_28,
    O => R1IN_2(46));
R1IN_2_ADD_1_CRY_29_Z7778: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_28,
    S => R1IN_2_ADD_1_AXB_29,
    LO => R1IN_2_ADD_1_CRY_29);
R1IN_2_ADD_1_S_28: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_28,
    CI => R1IN_2_ADD_1_CRY_27,
    O => R1IN_2(45));
R1IN_2_ADD_1_CRY_28_Z7780: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_27,
    S => R1IN_2_ADD_1_AXB_28,
    LO => R1IN_2_ADD_1_CRY_28);
R1IN_2_ADD_1_S_27: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_27,
    CI => R1IN_2_ADD_1_CRY_26,
    O => R1IN_2(44));
R1IN_2_ADD_1_CRY_27_Z7782: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_26,
    S => R1IN_2_ADD_1_AXB_27,
    LO => R1IN_2_ADD_1_CRY_27);
R1IN_2_ADD_1_S_26: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_26,
    CI => R1IN_2_ADD_1_CRY_25,
    O => R1IN_2(43));
R1IN_2_ADD_1_CRY_26_Z7784: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_25,
    S => R1IN_2_ADD_1_AXB_26,
    LO => R1IN_2_ADD_1_CRY_26);
R1IN_2_ADD_1_S_25: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_25,
    CI => R1IN_2_ADD_1_CRY_24,
    O => R1IN_2(42));
R1IN_2_ADD_1_CRY_25_Z7786: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_24,
    S => R1IN_2_ADD_1_AXB_25,
    LO => R1IN_2_ADD_1_CRY_25);
R1IN_2_ADD_1_S_24: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_24,
    CI => R1IN_2_ADD_1_CRY_23,
    O => R1IN_2(41));
R1IN_2_ADD_1_CRY_24_Z7788: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_23,
    S => R1IN_2_ADD_1_AXB_24,
    LO => R1IN_2_ADD_1_CRY_24);
R1IN_2_ADD_1_S_23: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_23,
    CI => R1IN_2_ADD_1_CRY_22,
    O => R1IN_2(40));
R1IN_2_ADD_1_CRY_23_Z7790: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_22,
    S => R1IN_2_ADD_1_AXB_23,
    LO => R1IN_2_ADD_1_CRY_23);
R1IN_2_ADD_1_S_22: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_22,
    CI => R1IN_2_ADD_1_CRY_21,
    O => R1IN_2(39));
R1IN_2_ADD_1_CRY_22_Z7792: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_21,
    S => R1IN_2_ADD_1_AXB_22,
    LO => R1IN_2_ADD_1_CRY_22);
R1IN_2_ADD_1_S_21: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_21,
    CI => R1IN_2_ADD_1_CRY_20,
    O => R1IN_2(38));
R1IN_2_ADD_1_CRY_21_Z7794: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_20,
    S => R1IN_2_ADD_1_AXB_21,
    LO => R1IN_2_ADD_1_CRY_21);
R1IN_2_ADD_1_S_20: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_20,
    CI => R1IN_2_ADD_1_CRY_19,
    O => R1IN_2(37));
R1IN_2_ADD_1_CRY_20_Z7796: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_19,
    S => R1IN_2_ADD_1_AXB_20,
    LO => R1IN_2_ADD_1_CRY_20);
R1IN_2_ADD_1_S_19: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_19,
    CI => R1IN_2_ADD_1_CRY_18,
    O => R1IN_2(36));
R1IN_2_ADD_1_CRY_19_Z7798: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_18,
    S => R1IN_2_ADD_1_AXB_19,
    LO => R1IN_2_ADD_1_CRY_19);
R1IN_2_ADD_1_S_18: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_18,
    CI => R1IN_2_ADD_1_CRY_17,
    O => R1IN_2(35));
R1IN_2_ADD_1_CRY_18_Z7800: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_17,
    S => R1IN_2_ADD_1_AXB_18,
    LO => R1IN_2_ADD_1_CRY_18);
R1IN_2_ADD_1_S_17: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_17,
    CI => R1IN_2_ADD_1_CRY_16,
    O => R1IN_2(34));
R1IN_2_ADD_1_CRY_17_Z7802: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_2_ADD_1_CRY_16,
    S => R1IN_2_ADD_1_AXB_17,
    LO => R1IN_2_ADD_1_CRY_17);
R1IN_2_ADD_1_S_16: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_16,
    CI => R1IN_2_ADD_1_CRY_15,
    O => R1IN_2(33));
R1IN_2_ADD_1_CRY_16_Z7804: MUXCY_L port map (
    DI => R1IN_2_2F(16),
    CI => R1IN_2_ADD_1_CRY_15,
    S => R1IN_2_ADD_1_AXB_16,
    LO => R1IN_2_ADD_1_CRY_16);
R1IN_2_ADD_1_S_15: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_15,
    CI => R1IN_2_ADD_1_CRY_14,
    O => R1IN_2(32));
R1IN_2_ADD_1_CRY_15_Z7806: MUXCY_L port map (
    DI => R1IN_2_2F(15),
    CI => R1IN_2_ADD_1_CRY_14,
    S => R1IN_2_ADD_1_AXB_15,
    LO => R1IN_2_ADD_1_CRY_15);
R1IN_2_ADD_1_S_14: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_14,
    CI => R1IN_2_ADD_1_CRY_13,
    O => R1IN_2(31));
R1IN_2_ADD_1_CRY_14_Z7808: MUXCY_L port map (
    DI => R1IN_2_2F(14),
    CI => R1IN_2_ADD_1_CRY_13,
    S => R1IN_2_ADD_1_AXB_14,
    LO => R1IN_2_ADD_1_CRY_14);
R1IN_2_ADD_1_S_13: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_13,
    CI => R1IN_2_ADD_1_CRY_12,
    O => R1IN_2(30));
R1IN_2_ADD_1_CRY_13_Z7810: MUXCY_L port map (
    DI => R1IN_2_2F(13),
    CI => R1IN_2_ADD_1_CRY_12,
    S => R1IN_2_ADD_1_AXB_13,
    LO => R1IN_2_ADD_1_CRY_13);
R1IN_2_ADD_1_S_12: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_12,
    CI => R1IN_2_ADD_1_CRY_11,
    O => R1IN_2(29));
R1IN_2_ADD_1_CRY_12_Z7812: MUXCY_L port map (
    DI => R1IN_2_2F(12),
    CI => R1IN_2_ADD_1_CRY_11,
    S => R1IN_2_ADD_1_AXB_12,
    LO => R1IN_2_ADD_1_CRY_12);
R1IN_2_ADD_1_S_11: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_11,
    CI => R1IN_2_ADD_1_CRY_10,
    O => R1IN_2(28));
R1IN_2_ADD_1_CRY_11_Z7814: MUXCY_L port map (
    DI => R1IN_2_2F(11),
    CI => R1IN_2_ADD_1_CRY_10,
    S => R1IN_2_ADD_1_AXB_11,
    LO => R1IN_2_ADD_1_CRY_11);
R1IN_2_ADD_1_S_10: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_10,
    CI => R1IN_2_ADD_1_CRY_9,
    O => R1IN_2(27));
R1IN_2_ADD_1_CRY_10_Z7816: MUXCY_L port map (
    DI => R1IN_2_2F(10),
    CI => R1IN_2_ADD_1_CRY_9,
    S => R1IN_2_ADD_1_AXB_10,
    LO => R1IN_2_ADD_1_CRY_10);
R1IN_2_ADD_1_S_9: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_9,
    CI => R1IN_2_ADD_1_CRY_8,
    O => R1IN_2(26));
R1IN_2_ADD_1_CRY_9_Z7818: MUXCY_L port map (
    DI => R1IN_2_2F(9),
    CI => R1IN_2_ADD_1_CRY_8,
    S => R1IN_2_ADD_1_AXB_9,
    LO => R1IN_2_ADD_1_CRY_9);
R1IN_2_ADD_1_S_8: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_8,
    CI => R1IN_2_ADD_1_CRY_7,
    O => R1IN_2(25));
R1IN_2_ADD_1_CRY_8_Z7820: MUXCY_L port map (
    DI => R1IN_2_2F(8),
    CI => R1IN_2_ADD_1_CRY_7,
    S => R1IN_2_ADD_1_AXB_8,
    LO => R1IN_2_ADD_1_CRY_8);
R1IN_2_ADD_1_S_7: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_7,
    CI => R1IN_2_ADD_1_CRY_6,
    O => R1IN_2(24));
R1IN_2_ADD_1_CRY_7_Z7822: MUXCY_L port map (
    DI => R1IN_2_2F(7),
    CI => R1IN_2_ADD_1_CRY_6,
    S => R1IN_2_ADD_1_AXB_7,
    LO => R1IN_2_ADD_1_CRY_7);
R1IN_2_ADD_1_S_6: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_6,
    CI => R1IN_2_ADD_1_CRY_5,
    O => R1IN_2(23));
R1IN_2_ADD_1_CRY_6_Z7824: MUXCY_L port map (
    DI => R1IN_2_2F(6),
    CI => R1IN_2_ADD_1_CRY_5,
    S => R1IN_2_ADD_1_AXB_6,
    LO => R1IN_2_ADD_1_CRY_6);
R1IN_2_ADD_1_S_5: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_5,
    CI => R1IN_2_ADD_1_CRY_4,
    O => R1IN_2(22));
R1IN_2_ADD_1_CRY_5_Z7826: MUXCY_L port map (
    DI => R1IN_2_2F(5),
    CI => R1IN_2_ADD_1_CRY_4,
    S => R1IN_2_ADD_1_AXB_5,
    LO => R1IN_2_ADD_1_CRY_5);
R1IN_2_ADD_1_S_4: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_4,
    CI => R1IN_2_ADD_1_CRY_3,
    O => R1IN_2(21));
R1IN_2_ADD_1_CRY_4_Z7828: MUXCY_L port map (
    DI => R1IN_2_2F(4),
    CI => R1IN_2_ADD_1_CRY_3,
    S => R1IN_2_ADD_1_AXB_4,
    LO => R1IN_2_ADD_1_CRY_4);
R1IN_2_ADD_1_S_3: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_3,
    CI => R1IN_2_ADD_1_CRY_2,
    O => R1IN_2(20));
R1IN_2_ADD_1_CRY_3_Z7830: MUXCY_L port map (
    DI => R1IN_2_2F(3),
    CI => R1IN_2_ADD_1_CRY_2,
    S => R1IN_2_ADD_1_AXB_3,
    LO => R1IN_2_ADD_1_CRY_3);
R1IN_2_ADD_1_S_2: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_2,
    CI => R1IN_2_ADD_1_CRY_1,
    O => R1IN_2(19));
R1IN_2_ADD_1_CRY_2_Z7832: MUXCY_L port map (
    DI => R1IN_2_2F(2),
    CI => R1IN_2_ADD_1_CRY_1,
    S => R1IN_2_ADD_1_AXB_2,
    LO => R1IN_2_ADD_1_CRY_2);
R1IN_2_ADD_1_S_1: XORCY port map (
    LI => R1IN_2_ADD_1_AXB_1,
    CI => R1IN_2_ADD_1_CRY_0,
    O => R1IN_2(18));
R1IN_2_ADD_1_CRY_1_Z7834: MUXCY_L port map (
    DI => R1IN_2_2F(1),
    CI => R1IN_2_ADD_1_CRY_0,
    S => R1IN_2_ADD_1_AXB_1,
    LO => R1IN_2_ADD_1_CRY_1);
R1IN_2_ADD_1_CRY_0_Z7835: MUXCY_L port map (
    DI => R1IN_2_ADD_1,
    CI => NN_1,
    S => R1IN_2(17),
    LO => R1IN_2_ADD_1_CRY_0);
R1IN_3_ADD_1_S_43: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_43,
    CI => R1IN_3_ADD_1_CRY_42,
    O => R1IN_3(60));
R1IN_3_ADD_1_S_42: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_42,
    CI => R1IN_3_ADD_1_CRY_41,
    O => R1IN_3(59));
R1IN_3_ADD_1_CRY_42_Z7838: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_41,
    S => R1IN_3_ADD_1_AXB_42,
    LO => R1IN_3_ADD_1_CRY_42);
R1IN_3_ADD_1_S_41: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_41,
    CI => R1IN_3_ADD_1_CRY_40,
    O => R1IN_3(58));
R1IN_3_ADD_1_CRY_41_Z7840: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_40,
    S => R1IN_3_ADD_1_AXB_41,
    LO => R1IN_3_ADD_1_CRY_41);
R1IN_3_ADD_1_S_40: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_40,
    CI => R1IN_3_ADD_1_CRY_39,
    O => R1IN_3(57));
R1IN_3_ADD_1_CRY_40_Z7842: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_39,
    S => R1IN_3_ADD_1_AXB_40,
    LO => R1IN_3_ADD_1_CRY_40);
R1IN_3_ADD_1_S_39: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_39,
    CI => R1IN_3_ADD_1_CRY_38,
    O => R1IN_3(56));
R1IN_3_ADD_1_CRY_39_Z7844: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_38,
    S => R1IN_3_ADD_1_AXB_39,
    LO => R1IN_3_ADD_1_CRY_39);
R1IN_3_ADD_1_S_38: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_38,
    CI => R1IN_3_ADD_1_CRY_37,
    O => R1IN_3(55));
R1IN_3_ADD_1_CRY_38_Z7846: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_37,
    S => R1IN_3_ADD_1_AXB_38,
    LO => R1IN_3_ADD_1_CRY_38);
R1IN_3_ADD_1_S_37: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_37,
    CI => R1IN_3_ADD_1_CRY_36,
    O => R1IN_3(54));
R1IN_3_ADD_1_CRY_37_Z7848: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_36,
    S => R1IN_3_ADD_1_AXB_37,
    LO => R1IN_3_ADD_1_CRY_37);
R1IN_3_ADD_1_S_36: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_36,
    CI => R1IN_3_ADD_1_CRY_35,
    O => R1IN_3(53));
R1IN_3_ADD_1_CRY_36_Z7850: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_35,
    S => R1IN_3_ADD_1_AXB_36,
    LO => R1IN_3_ADD_1_CRY_36);
R1IN_3_ADD_1_S_35: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_35,
    CI => R1IN_3_ADD_1_CRY_34,
    O => R1IN_3(52));
R1IN_3_ADD_1_CRY_35_Z7852: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_34,
    S => R1IN_3_ADD_1_AXB_35,
    LO => R1IN_3_ADD_1_CRY_35);
R1IN_3_ADD_1_S_34: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_34,
    CI => R1IN_3_ADD_1_CRY_33,
    O => R1IN_3(51));
R1IN_3_ADD_1_CRY_34_Z7854: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_33,
    S => R1IN_3_ADD_1_AXB_34,
    LO => R1IN_3_ADD_1_CRY_34);
R1IN_3_ADD_1_S_33: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_33,
    CI => R1IN_3_ADD_1_CRY_32,
    O => R1IN_3(50));
R1IN_3_ADD_1_CRY_33_Z7856: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_32,
    S => R1IN_3_ADD_1_AXB_33,
    LO => R1IN_3_ADD_1_CRY_33);
R1IN_3_ADD_1_S_32: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_32,
    CI => R1IN_3_ADD_1_CRY_31,
    O => R1IN_3(49));
R1IN_3_ADD_1_CRY_32_Z7858: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_31,
    S => R1IN_3_ADD_1_AXB_32,
    LO => R1IN_3_ADD_1_CRY_32);
R1IN_3_ADD_1_S_31: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_31,
    CI => R1IN_3_ADD_1_CRY_30,
    O => R1IN_3(48));
R1IN_3_ADD_1_CRY_31_Z7860: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_30,
    S => R1IN_3_ADD_1_AXB_31,
    LO => R1IN_3_ADD_1_CRY_31);
R1IN_3_ADD_1_S_30: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_30,
    CI => R1IN_3_ADD_1_CRY_29,
    O => R1IN_3(47));
R1IN_3_ADD_1_CRY_30_Z7862: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_29,
    S => R1IN_3_ADD_1_AXB_30,
    LO => R1IN_3_ADD_1_CRY_30);
R1IN_3_ADD_1_S_29: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_29,
    CI => R1IN_3_ADD_1_CRY_28,
    O => R1IN_3(46));
R1IN_3_ADD_1_CRY_29_Z7864: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_28,
    S => R1IN_3_ADD_1_AXB_29,
    LO => R1IN_3_ADD_1_CRY_29);
R1IN_3_ADD_1_S_28: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_28,
    CI => R1IN_3_ADD_1_CRY_27,
    O => R1IN_3(45));
R1IN_3_ADD_1_CRY_28_Z7866: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_27,
    S => R1IN_3_ADD_1_AXB_28,
    LO => R1IN_3_ADD_1_CRY_28);
R1IN_3_ADD_1_S_27: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_27,
    CI => R1IN_3_ADD_1_CRY_26,
    O => R1IN_3(44));
R1IN_3_ADD_1_CRY_27_Z7868: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_26,
    S => R1IN_3_ADD_1_AXB_27,
    LO => R1IN_3_ADD_1_CRY_27);
R1IN_3_ADD_1_S_26: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_26,
    CI => R1IN_3_ADD_1_CRY_25,
    O => R1IN_3(43));
R1IN_3_ADD_1_CRY_26_Z7870: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_25,
    S => R1IN_3_ADD_1_AXB_26,
    LO => R1IN_3_ADD_1_CRY_26);
R1IN_3_ADD_1_S_25: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_25,
    CI => R1IN_3_ADD_1_CRY_24,
    O => R1IN_3(42));
R1IN_3_ADD_1_CRY_25_Z7872: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_24,
    S => R1IN_3_ADD_1_AXB_25,
    LO => R1IN_3_ADD_1_CRY_25);
R1IN_3_ADD_1_S_24: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_24,
    CI => R1IN_3_ADD_1_CRY_23,
    O => R1IN_3(41));
R1IN_3_ADD_1_CRY_24_Z7874: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_23,
    S => R1IN_3_ADD_1_AXB_24,
    LO => R1IN_3_ADD_1_CRY_24);
R1IN_3_ADD_1_S_23: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_23,
    CI => R1IN_3_ADD_1_CRY_22,
    O => R1IN_3(40));
R1IN_3_ADD_1_CRY_23_Z7876: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_22,
    S => R1IN_3_ADD_1_AXB_23,
    LO => R1IN_3_ADD_1_CRY_23);
R1IN_3_ADD_1_S_22: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_22,
    CI => R1IN_3_ADD_1_CRY_21,
    O => R1IN_3(39));
R1IN_3_ADD_1_CRY_22_Z7878: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_21,
    S => R1IN_3_ADD_1_AXB_22,
    LO => R1IN_3_ADD_1_CRY_22);
R1IN_3_ADD_1_S_21: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_21,
    CI => R1IN_3_ADD_1_CRY_20,
    O => R1IN_3(38));
R1IN_3_ADD_1_CRY_21_Z7880: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_20,
    S => R1IN_3_ADD_1_AXB_21,
    LO => R1IN_3_ADD_1_CRY_21);
R1IN_3_ADD_1_S_20: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_20,
    CI => R1IN_3_ADD_1_CRY_19,
    O => R1IN_3(37));
R1IN_3_ADD_1_CRY_20_Z7882: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_19,
    S => R1IN_3_ADD_1_AXB_20,
    LO => R1IN_3_ADD_1_CRY_20);
R1IN_3_ADD_1_S_19: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_19,
    CI => R1IN_3_ADD_1_CRY_18,
    O => R1IN_3(36));
R1IN_3_ADD_1_CRY_19_Z7884: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_18,
    S => R1IN_3_ADD_1_AXB_19,
    LO => R1IN_3_ADD_1_CRY_19);
R1IN_3_ADD_1_S_18: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_18,
    CI => R1IN_3_ADD_1_CRY_17,
    O => R1IN_3(35));
R1IN_3_ADD_1_CRY_18_Z7886: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_17,
    S => R1IN_3_ADD_1_AXB_18,
    LO => R1IN_3_ADD_1_CRY_18);
R1IN_3_ADD_1_S_17: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_17,
    CI => R1IN_3_ADD_1_CRY_16,
    O => R1IN_3(34));
R1IN_3_ADD_1_CRY_17_Z7888: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_3_ADD_1_CRY_16,
    S => R1IN_3_ADD_1_AXB_17,
    LO => R1IN_3_ADD_1_CRY_17);
R1IN_3_ADD_1_S_16: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_16,
    CI => R1IN_3_ADD_1_CRY_15,
    O => R1IN_3(33));
R1IN_3_ADD_1_CRY_16_Z7890: MUXCY_L port map (
    DI => R1IN_3_2F(16),
    CI => R1IN_3_ADD_1_CRY_15,
    S => R1IN_3_ADD_1_AXB_16,
    LO => R1IN_3_ADD_1_CRY_16);
R1IN_3_ADD_1_S_15: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_15,
    CI => R1IN_3_ADD_1_CRY_14,
    O => R1IN_3(32));
R1IN_3_ADD_1_CRY_15_Z7892: MUXCY_L port map (
    DI => R1IN_3_2F(15),
    CI => R1IN_3_ADD_1_CRY_14,
    S => R1IN_3_ADD_1_AXB_15,
    LO => R1IN_3_ADD_1_CRY_15);
R1IN_3_ADD_1_S_14: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_14,
    CI => R1IN_3_ADD_1_CRY_13,
    O => R1IN_3(31));
R1IN_3_ADD_1_CRY_14_Z7894: MUXCY_L port map (
    DI => R1IN_3_2F(14),
    CI => R1IN_3_ADD_1_CRY_13,
    S => R1IN_3_ADD_1_AXB_14,
    LO => R1IN_3_ADD_1_CRY_14);
R1IN_3_ADD_1_S_13: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_13,
    CI => R1IN_3_ADD_1_CRY_12,
    O => R1IN_3(30));
R1IN_3_ADD_1_CRY_13_Z7896: MUXCY_L port map (
    DI => R1IN_3_2F(13),
    CI => R1IN_3_ADD_1_CRY_12,
    S => R1IN_3_ADD_1_AXB_13,
    LO => R1IN_3_ADD_1_CRY_13);
R1IN_3_ADD_1_S_12: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_12,
    CI => R1IN_3_ADD_1_CRY_11,
    O => R1IN_3(29));
R1IN_3_ADD_1_CRY_12_Z7898: MUXCY_L port map (
    DI => R1IN_3_2F(12),
    CI => R1IN_3_ADD_1_CRY_11,
    S => R1IN_3_ADD_1_AXB_12,
    LO => R1IN_3_ADD_1_CRY_12);
R1IN_3_ADD_1_S_11: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_11,
    CI => R1IN_3_ADD_1_CRY_10,
    O => R1IN_3(28));
R1IN_3_ADD_1_CRY_11_Z7900: MUXCY_L port map (
    DI => R1IN_3_2F(11),
    CI => R1IN_3_ADD_1_CRY_10,
    S => R1IN_3_ADD_1_AXB_11,
    LO => R1IN_3_ADD_1_CRY_11);
R1IN_3_ADD_1_S_10: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_10,
    CI => R1IN_3_ADD_1_CRY_9,
    O => R1IN_3(27));
R1IN_3_ADD_1_CRY_10_Z7902: MUXCY_L port map (
    DI => R1IN_3_2F(10),
    CI => R1IN_3_ADD_1_CRY_9,
    S => R1IN_3_ADD_1_AXB_10,
    LO => R1IN_3_ADD_1_CRY_10);
R1IN_3_ADD_1_S_9: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_9,
    CI => R1IN_3_ADD_1_CRY_8,
    O => R1IN_3(26));
R1IN_3_ADD_1_CRY_9_Z7904: MUXCY_L port map (
    DI => R1IN_3_2F(9),
    CI => R1IN_3_ADD_1_CRY_8,
    S => R1IN_3_ADD_1_AXB_9,
    LO => R1IN_3_ADD_1_CRY_9);
R1IN_3_ADD_1_S_8: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_8,
    CI => R1IN_3_ADD_1_CRY_7,
    O => R1IN_3(25));
R1IN_3_ADD_1_CRY_8_Z7906: MUXCY_L port map (
    DI => R1IN_3_2F(8),
    CI => R1IN_3_ADD_1_CRY_7,
    S => R1IN_3_ADD_1_AXB_8,
    LO => R1IN_3_ADD_1_CRY_8);
R1IN_3_ADD_1_S_7: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_7,
    CI => R1IN_3_ADD_1_CRY_6,
    O => R1IN_3(24));
R1IN_3_ADD_1_CRY_7_Z7908: MUXCY_L port map (
    DI => R1IN_3_2F(7),
    CI => R1IN_3_ADD_1_CRY_6,
    S => R1IN_3_ADD_1_AXB_7,
    LO => R1IN_3_ADD_1_CRY_7);
R1IN_3_ADD_1_S_6: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_6,
    CI => R1IN_3_ADD_1_CRY_5,
    O => R1IN_3(23));
R1IN_3_ADD_1_CRY_6_Z7910: MUXCY_L port map (
    DI => R1IN_3_2F(6),
    CI => R1IN_3_ADD_1_CRY_5,
    S => R1IN_3_ADD_1_AXB_6,
    LO => R1IN_3_ADD_1_CRY_6);
R1IN_3_ADD_1_S_5: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_5,
    CI => R1IN_3_ADD_1_CRY_4,
    O => R1IN_3(22));
R1IN_3_ADD_1_CRY_5_Z7912: MUXCY_L port map (
    DI => R1IN_3_2F(5),
    CI => R1IN_3_ADD_1_CRY_4,
    S => R1IN_3_ADD_1_AXB_5,
    LO => R1IN_3_ADD_1_CRY_5);
R1IN_3_ADD_1_S_4: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_4,
    CI => R1IN_3_ADD_1_CRY_3,
    O => R1IN_3(21));
R1IN_3_ADD_1_CRY_4_Z7914: MUXCY_L port map (
    DI => R1IN_3_2F(4),
    CI => R1IN_3_ADD_1_CRY_3,
    S => R1IN_3_ADD_1_AXB_4,
    LO => R1IN_3_ADD_1_CRY_4);
R1IN_3_ADD_1_S_3: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_3,
    CI => R1IN_3_ADD_1_CRY_2,
    O => R1IN_3(20));
R1IN_3_ADD_1_CRY_3_Z7916: MUXCY_L port map (
    DI => R1IN_3_2F(3),
    CI => R1IN_3_ADD_1_CRY_2,
    S => R1IN_3_ADD_1_AXB_3,
    LO => R1IN_3_ADD_1_CRY_3);
R1IN_3_ADD_1_S_2: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_2,
    CI => R1IN_3_ADD_1_CRY_1,
    O => R1IN_3(19));
R1IN_3_ADD_1_CRY_2_Z7918: MUXCY_L port map (
    DI => R1IN_3_2F(2),
    CI => R1IN_3_ADD_1_CRY_1,
    S => R1IN_3_ADD_1_AXB_2,
    LO => R1IN_3_ADD_1_CRY_2);
R1IN_3_ADD_1_S_1: XORCY port map (
    LI => R1IN_3_ADD_1_AXB_1,
    CI => R1IN_3_ADD_1_CRY_0,
    O => R1IN_3(18));
R1IN_3_ADD_1_CRY_1_Z7920: MUXCY_L port map (
    DI => R1IN_3_2F(1),
    CI => R1IN_3_ADD_1_CRY_0,
    S => R1IN_3_ADD_1_AXB_1,
    LO => R1IN_3_ADD_1_CRY_1);
R1IN_3_ADD_1_CRY_0_Z7921: MUXCY_L port map (
    DI => R1IN_3_ADD_1,
    CI => NN_1,
    S => R1IN_3(17),
    LO => R1IN_3_ADD_1_CRY_0);
R1IN_ADD_1_1_0_S_28_Z7922: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_28,
    CI => R1IN_ADD_1_1_0_CRY_27,
    O => R1IN_ADD_1_1_0_S_28);
R1IN_ADD_1_1_0_CRY_28_Z7923: MUXCY port map (
    DI => R1IN_3(60),
    CI => R1IN_ADD_1_1_0_CRY_27,
    S => R1IN_ADD_1_1_0_AXB_28,
    O => R1IN_ADD_1_1_0_CRY_28);
R1IN_ADD_1_1_0_S_27_Z7924: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_27,
    CI => R1IN_ADD_1_1_0_CRY_26,
    O => R1IN_ADD_1_1_0_S_27);
R1IN_ADD_1_1_0_CRY_27_Z7925: MUXCY_L port map (
    DI => R1IN_3(59),
    CI => R1IN_ADD_1_1_0_CRY_26,
    S => R1IN_ADD_1_1_0_AXB_27,
    LO => R1IN_ADD_1_1_0_CRY_27);
R1IN_ADD_1_1_0_S_26_Z7926: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_26,
    CI => R1IN_ADD_1_1_0_CRY_25,
    O => R1IN_ADD_1_1_0_S_26);
R1IN_ADD_1_1_0_CRY_26_Z7927: MUXCY_L port map (
    DI => R1IN_3(58),
    CI => R1IN_ADD_1_1_0_CRY_25,
    S => R1IN_ADD_1_1_0_AXB_26,
    LO => R1IN_ADD_1_1_0_CRY_26);
R1IN_ADD_1_1_0_S_25_Z7928: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_25,
    CI => R1IN_ADD_1_1_0_CRY_24,
    O => R1IN_ADD_1_1_0_S_25);
R1IN_ADD_1_1_0_CRY_25_Z7929: MUXCY_L port map (
    DI => R1IN_3(57),
    CI => R1IN_ADD_1_1_0_CRY_24,
    S => R1IN_ADD_1_1_0_AXB_25,
    LO => R1IN_ADD_1_1_0_CRY_25);
R1IN_ADD_1_1_0_S_24_Z7930: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_24,
    CI => R1IN_ADD_1_1_0_CRY_23,
    O => R1IN_ADD_1_1_0_S_24);
R1IN_ADD_1_1_0_CRY_24_Z7931: MUXCY_L port map (
    DI => R1IN_3(56),
    CI => R1IN_ADD_1_1_0_CRY_23,
    S => R1IN_ADD_1_1_0_AXB_24,
    LO => R1IN_ADD_1_1_0_CRY_24);
R1IN_ADD_1_1_0_S_23_Z7932: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_23,
    CI => R1IN_ADD_1_1_0_CRY_22,
    O => R1IN_ADD_1_1_0_S_23);
R1IN_ADD_1_1_0_CRY_23_Z7933: MUXCY_L port map (
    DI => R1IN_3(55),
    CI => R1IN_ADD_1_1_0_CRY_22,
    S => R1IN_ADD_1_1_0_AXB_23,
    LO => R1IN_ADD_1_1_0_CRY_23);
R1IN_ADD_1_1_0_S_22_Z7934: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_22,
    CI => R1IN_ADD_1_1_0_CRY_21,
    O => R1IN_ADD_1_1_0_S_22);
R1IN_ADD_1_1_0_CRY_22_Z7935: MUXCY_L port map (
    DI => R1IN_3(54),
    CI => R1IN_ADD_1_1_0_CRY_21,
    S => R1IN_ADD_1_1_0_AXB_22,
    LO => R1IN_ADD_1_1_0_CRY_22);
R1IN_ADD_1_1_0_S_21_Z7936: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_21,
    CI => R1IN_ADD_1_1_0_CRY_20,
    O => R1IN_ADD_1_1_0_S_21);
R1IN_ADD_1_1_0_CRY_21_Z7937: MUXCY_L port map (
    DI => R1IN_3(53),
    CI => R1IN_ADD_1_1_0_CRY_20,
    S => R1IN_ADD_1_1_0_AXB_21,
    LO => R1IN_ADD_1_1_0_CRY_21);
R1IN_ADD_1_1_0_S_20: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_20,
    CI => R1IN_ADD_1_1_0_CRY_19,
    O => N_1913);
R1IN_ADD_1_1_0_CRY_20_Z7939: MUXCY_L port map (
    DI => R1IN_3(52),
    CI => R1IN_ADD_1_1_0_CRY_19,
    S => R1IN_ADD_1_1_0_AXB_20,
    LO => R1IN_ADD_1_1_0_CRY_20);
R1IN_ADD_1_1_0_S_19: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_19,
    CI => R1IN_ADD_1_1_0_CRY_18,
    O => N_1912);
R1IN_ADD_1_1_0_CRY_19_Z7941: MUXCY_L port map (
    DI => R1IN_3(51),
    CI => R1IN_ADD_1_1_0_CRY_18,
    S => R1IN_ADD_1_1_0_AXB_19,
    LO => R1IN_ADD_1_1_0_CRY_19);
R1IN_ADD_1_1_0_S_18: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_18,
    CI => R1IN_ADD_1_1_0_CRY_17,
    O => N_1911);
R1IN_ADD_1_1_0_CRY_18_Z7943: MUXCY_L port map (
    DI => R1IN_3(50),
    CI => R1IN_ADD_1_1_0_CRY_17,
    S => R1IN_ADD_1_1_0_AXB_18,
    LO => R1IN_ADD_1_1_0_CRY_18);
R1IN_ADD_1_1_0_S_17: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_17,
    CI => R1IN_ADD_1_1_0_CRY_16,
    O => N_1910);
R1IN_ADD_1_1_0_CRY_17_Z7945: MUXCY_L port map (
    DI => R1IN_3(49),
    CI => R1IN_ADD_1_1_0_CRY_16,
    S => R1IN_ADD_1_1_0_AXB_17,
    LO => R1IN_ADD_1_1_0_CRY_17);
R1IN_ADD_1_1_0_S_16: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_16,
    CI => R1IN_ADD_1_1_0_CRY_15,
    O => N_1909);
R1IN_ADD_1_1_0_CRY_16_Z7947: MUXCY_L port map (
    DI => R1IN_3(48),
    CI => R1IN_ADD_1_1_0_CRY_15,
    S => R1IN_ADD_1_1_0_AXB_16,
    LO => R1IN_ADD_1_1_0_CRY_16);
R1IN_ADD_1_1_0_S_15: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_15,
    CI => R1IN_ADD_1_1_0_CRY_14,
    O => N_1908);
R1IN_ADD_1_1_0_CRY_15_Z7949: MUXCY_L port map (
    DI => R1IN_3(47),
    CI => R1IN_ADD_1_1_0_CRY_14,
    S => R1IN_ADD_1_1_0_AXB_15,
    LO => R1IN_ADD_1_1_0_CRY_15);
R1IN_ADD_1_1_0_S_14: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_14,
    CI => R1IN_ADD_1_1_0_CRY_13,
    O => N_1907);
R1IN_ADD_1_1_0_CRY_14_Z7951: MUXCY_L port map (
    DI => R1IN_3(46),
    CI => R1IN_ADD_1_1_0_CRY_13,
    S => R1IN_ADD_1_1_0_AXB_14,
    LO => R1IN_ADD_1_1_0_CRY_14);
R1IN_ADD_1_1_0_S_13: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_13,
    CI => R1IN_ADD_1_1_0_CRY_12,
    O => N_1906);
R1IN_ADD_1_1_0_CRY_13_Z7953: MUXCY_L port map (
    DI => R1IN_3(45),
    CI => R1IN_ADD_1_1_0_CRY_12,
    S => R1IN_ADD_1_1_0_AXB_13,
    LO => R1IN_ADD_1_1_0_CRY_13);
R1IN_ADD_1_1_0_S_12: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_12,
    CI => R1IN_ADD_1_1_0_CRY_11,
    O => N_1905);
R1IN_ADD_1_1_0_CRY_12_Z7955: MUXCY_L port map (
    DI => R1IN_3(44),
    CI => R1IN_ADD_1_1_0_CRY_11,
    S => R1IN_ADD_1_1_0_AXB_12,
    LO => R1IN_ADD_1_1_0_CRY_12);
R1IN_ADD_1_1_0_S_11: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_11,
    CI => R1IN_ADD_1_1_0_CRY_10,
    O => N_1904);
R1IN_ADD_1_1_0_CRY_11_Z7957: MUXCY_L port map (
    DI => R1IN_3(43),
    CI => R1IN_ADD_1_1_0_CRY_10,
    S => R1IN_ADD_1_1_0_AXB_11,
    LO => R1IN_ADD_1_1_0_CRY_11);
R1IN_ADD_1_1_0_S_10: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_10,
    CI => R1IN_ADD_1_1_0_CRY_9,
    O => N_1903);
R1IN_ADD_1_1_0_CRY_10_Z7959: MUXCY_L port map (
    DI => R1IN_3(42),
    CI => R1IN_ADD_1_1_0_CRY_9,
    S => R1IN_ADD_1_1_0_AXB_10,
    LO => R1IN_ADD_1_1_0_CRY_10);
R1IN_ADD_1_1_0_S_9: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_9,
    CI => R1IN_ADD_1_1_0_CRY_8,
    O => N_1902);
R1IN_ADD_1_1_0_CRY_9_Z7961: MUXCY_L port map (
    DI => R1IN_3(41),
    CI => R1IN_ADD_1_1_0_CRY_8,
    S => R1IN_ADD_1_1_0_AXB_9,
    LO => R1IN_ADD_1_1_0_CRY_9);
R1IN_ADD_1_1_0_S_8: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_8,
    CI => R1IN_ADD_1_1_0_CRY_7,
    O => N_1901);
R1IN_ADD_1_1_0_CRY_8_Z7963: MUXCY_L port map (
    DI => R1IN_3(40),
    CI => R1IN_ADD_1_1_0_CRY_7,
    S => R1IN_ADD_1_1_0_AXB_8,
    LO => R1IN_ADD_1_1_0_CRY_8);
R1IN_ADD_1_1_0_S_7: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_7,
    CI => R1IN_ADD_1_1_0_CRY_6,
    O => N_1900);
R1IN_ADD_1_1_0_CRY_7_Z7965: MUXCY_L port map (
    DI => R1IN_3(39),
    CI => R1IN_ADD_1_1_0_CRY_6,
    S => R1IN_ADD_1_1_0_AXB_7,
    LO => R1IN_ADD_1_1_0_CRY_7);
R1IN_ADD_1_1_0_S_6: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_6,
    CI => R1IN_ADD_1_1_0_CRY_5,
    O => N_1899);
R1IN_ADD_1_1_0_CRY_6_Z7967: MUXCY_L port map (
    DI => R1IN_3(38),
    CI => R1IN_ADD_1_1_0_CRY_5,
    S => R1IN_ADD_1_1_0_AXB_6,
    LO => R1IN_ADD_1_1_0_CRY_6);
R1IN_ADD_1_1_0_S_5: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_5,
    CI => R1IN_ADD_1_1_0_CRY_4,
    O => N_1898);
R1IN_ADD_1_1_0_CRY_5_Z7969: MUXCY_L port map (
    DI => R1IN_3(37),
    CI => R1IN_ADD_1_1_0_CRY_4,
    S => R1IN_ADD_1_1_0_AXB_5,
    LO => R1IN_ADD_1_1_0_CRY_5);
R1IN_ADD_1_1_0_S_4: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_4,
    CI => R1IN_ADD_1_1_0_CRY_3,
    O => N_1897);
R1IN_ADD_1_1_0_CRY_4_Z7971: MUXCY_L port map (
    DI => R1IN_3(36),
    CI => R1IN_ADD_1_1_0_CRY_3,
    S => R1IN_ADD_1_1_0_AXB_4,
    LO => R1IN_ADD_1_1_0_CRY_4);
R1IN_ADD_1_1_0_S_3: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_3,
    CI => R1IN_ADD_1_1_0_CRY_2,
    O => N_1896);
R1IN_ADD_1_1_0_CRY_3_Z7973: MUXCY_L port map (
    DI => R1IN_3(35),
    CI => R1IN_ADD_1_1_0_CRY_2,
    S => R1IN_ADD_1_1_0_AXB_3,
    LO => R1IN_ADD_1_1_0_CRY_3);
R1IN_ADD_1_1_0_S_2: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_2,
    CI => R1IN_ADD_1_1_0_CRY_1,
    O => N_1895);
R1IN_ADD_1_1_0_CRY_2_Z7975: MUXCY_L port map (
    DI => R1IN_3(34),
    CI => R1IN_ADD_1_1_0_CRY_1,
    S => R1IN_ADD_1_1_0_AXB_2,
    LO => R1IN_ADD_1_1_0_CRY_2);
R1IN_ADD_1_1_0_S_1: XORCY port map (
    LI => R1IN_ADD_1_1_0_AXB_1,
    CI => R1IN_ADD_1_1_0_CRY_0,
    O => N_1894);
R1IN_ADD_1_1_0_CRY_1_Z7977: MUXCY_L port map (
    DI => R1IN_3(33),
    CI => R1IN_ADD_1_1_0_CRY_0,
    S => R1IN_ADD_1_1_0_AXB_1,
    LO => R1IN_ADD_1_1_0_CRY_1);
R1IN_ADD_1_1_0_CRY_0_Z7978: MUXCY_L port map (
    DI => R1IN_3(32),
    CI => NN_2,
    S => R1IN_ADD_1_1_0_AXB_0,
    LO => R1IN_ADD_1_1_0_CRY_0);
R1IN_ADD_1_1_S_28_Z7979: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_28,
    CI => R1IN_ADD_1_1_CRY_27,
    O => R1IN_ADD_1_1_S_28);
R1IN_ADD_1_1_S_27_Z7980: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_27,
    CI => R1IN_ADD_1_1_CRY_26,
    O => R1IN_ADD_1_1_S_27);
R1IN_ADD_1_1_CRY_27_Z7981: MUXCY_L port map (
    DI => R1IN_3(59),
    CI => R1IN_ADD_1_1_CRY_26,
    S => R1IN_ADD_1_1_AXB_27,
    LO => R1IN_ADD_1_1_CRY_27);
R1IN_ADD_1_1_S_26_Z7982: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_26,
    CI => R1IN_ADD_1_1_CRY_25,
    O => R1IN_ADD_1_1_S_26);
R1IN_ADD_1_1_CRY_26_Z7983: MUXCY_L port map (
    DI => R1IN_3(58),
    CI => R1IN_ADD_1_1_CRY_25,
    S => R1IN_ADD_1_1_AXB_26,
    LO => R1IN_ADD_1_1_CRY_26);
R1IN_ADD_1_1_S_25_Z7984: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_25,
    CI => R1IN_ADD_1_1_CRY_24,
    O => R1IN_ADD_1_1_S_25);
R1IN_ADD_1_1_CRY_25_Z7985: MUXCY_L port map (
    DI => R1IN_3(57),
    CI => R1IN_ADD_1_1_CRY_24,
    S => R1IN_ADD_1_1_AXB_25,
    LO => R1IN_ADD_1_1_CRY_25);
R1IN_ADD_1_1_S_24_Z7986: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_24,
    CI => R1IN_ADD_1_1_CRY_23,
    O => R1IN_ADD_1_1_S_24);
R1IN_ADD_1_1_CRY_24_Z7987: MUXCY_L port map (
    DI => R1IN_3(56),
    CI => R1IN_ADD_1_1_CRY_23,
    S => R1IN_ADD_1_1_AXB_24,
    LO => R1IN_ADD_1_1_CRY_24);
R1IN_ADD_1_1_S_23_Z7988: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_23,
    CI => R1IN_ADD_1_1_CRY_22,
    O => R1IN_ADD_1_1_S_23);
R1IN_ADD_1_1_CRY_23_Z7989: MUXCY_L port map (
    DI => R1IN_3(55),
    CI => R1IN_ADD_1_1_CRY_22,
    S => R1IN_ADD_1_1_AXB_23,
    LO => R1IN_ADD_1_1_CRY_23);
R1IN_ADD_1_1_S_22_Z7990: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_22,
    CI => R1IN_ADD_1_1_CRY_21,
    O => R1IN_ADD_1_1_S_22);
R1IN_ADD_1_1_CRY_22_Z7991: MUXCY_L port map (
    DI => R1IN_3(54),
    CI => R1IN_ADD_1_1_CRY_21,
    S => R1IN_ADD_1_1_AXB_22,
    LO => R1IN_ADD_1_1_CRY_22);
R1IN_ADD_1_1_S_21_Z7992: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_21,
    CI => R1IN_ADD_1_1_CRY_20,
    O => R1IN_ADD_1_1_S_21);
R1IN_ADD_1_1_CRY_21_Z7993: MUXCY_L port map (
    DI => R1IN_3(53),
    CI => R1IN_ADD_1_1_CRY_20,
    S => R1IN_ADD_1_1_AXB_21,
    LO => R1IN_ADD_1_1_CRY_21);
R1IN_ADD_1_1_S_20: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_20,
    CI => R1IN_ADD_1_1_CRY_19,
    O => N_1577);
R1IN_ADD_1_1_CRY_20_Z7995: MUXCY_L port map (
    DI => R1IN_3(52),
    CI => R1IN_ADD_1_1_CRY_19,
    S => R1IN_ADD_1_1_AXB_20,
    LO => R1IN_ADD_1_1_CRY_20);
R1IN_ADD_1_1_S_19: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_19,
    CI => R1IN_ADD_1_1_CRY_18,
    O => N_1575);
R1IN_ADD_1_1_CRY_19_Z7997: MUXCY_L port map (
    DI => R1IN_3(51),
    CI => R1IN_ADD_1_1_CRY_18,
    S => R1IN_ADD_1_1_AXB_19,
    LO => R1IN_ADD_1_1_CRY_19);
R1IN_ADD_1_1_S_18: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_18,
    CI => R1IN_ADD_1_1_CRY_17,
    O => N_1573);
R1IN_ADD_1_1_CRY_18_Z7999: MUXCY_L port map (
    DI => R1IN_3(50),
    CI => R1IN_ADD_1_1_CRY_17,
    S => R1IN_ADD_1_1_AXB_18,
    LO => R1IN_ADD_1_1_CRY_18);
R1IN_ADD_1_1_S_17: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_17,
    CI => R1IN_ADD_1_1_CRY_16,
    O => N_1571);
R1IN_ADD_1_1_CRY_17_Z8001: MUXCY_L port map (
    DI => R1IN_3(49),
    CI => R1IN_ADD_1_1_CRY_16,
    S => R1IN_ADD_1_1_AXB_17,
    LO => R1IN_ADD_1_1_CRY_17);
R1IN_ADD_1_1_S_16: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_16,
    CI => R1IN_ADD_1_1_CRY_15,
    O => N_1569);
R1IN_ADD_1_1_CRY_16_Z8003: MUXCY_L port map (
    DI => R1IN_3(48),
    CI => R1IN_ADD_1_1_CRY_15,
    S => R1IN_ADD_1_1_AXB_16,
    LO => R1IN_ADD_1_1_CRY_16);
R1IN_ADD_1_1_S_15: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_15,
    CI => R1IN_ADD_1_1_CRY_14,
    O => N_1567);
R1IN_ADD_1_1_CRY_15_Z8005: MUXCY_L port map (
    DI => R1IN_3(47),
    CI => R1IN_ADD_1_1_CRY_14,
    S => R1IN_ADD_1_1_AXB_15,
    LO => R1IN_ADD_1_1_CRY_15);
R1IN_ADD_1_1_S_14: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_14,
    CI => R1IN_ADD_1_1_CRY_13,
    O => N_1565);
R1IN_ADD_1_1_CRY_14_Z8007: MUXCY_L port map (
    DI => R1IN_3(46),
    CI => R1IN_ADD_1_1_CRY_13,
    S => R1IN_ADD_1_1_AXB_14,
    LO => R1IN_ADD_1_1_CRY_14);
R1IN_ADD_1_1_S_13: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_13,
    CI => R1IN_ADD_1_1_CRY_12,
    O => N_1563);
R1IN_ADD_1_1_CRY_13_Z8009: MUXCY_L port map (
    DI => R1IN_3(45),
    CI => R1IN_ADD_1_1_CRY_12,
    S => R1IN_ADD_1_1_AXB_13,
    LO => R1IN_ADD_1_1_CRY_13);
R1IN_ADD_1_1_S_12: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_12,
    CI => R1IN_ADD_1_1_CRY_11,
    O => N_1561);
R1IN_ADD_1_1_CRY_12_Z8011: MUXCY_L port map (
    DI => R1IN_3(44),
    CI => R1IN_ADD_1_1_CRY_11,
    S => R1IN_ADD_1_1_AXB_12,
    LO => R1IN_ADD_1_1_CRY_12);
R1IN_ADD_1_1_S_11: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_11,
    CI => R1IN_ADD_1_1_CRY_10,
    O => N_1559);
R1IN_ADD_1_1_CRY_11_Z8013: MUXCY_L port map (
    DI => R1IN_3(43),
    CI => R1IN_ADD_1_1_CRY_10,
    S => R1IN_ADD_1_1_AXB_11,
    LO => R1IN_ADD_1_1_CRY_11);
R1IN_ADD_1_1_S_10: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_10,
    CI => R1IN_ADD_1_1_CRY_9,
    O => N_1557);
R1IN_ADD_1_1_CRY_10_Z8015: MUXCY_L port map (
    DI => R1IN_3(42),
    CI => R1IN_ADD_1_1_CRY_9,
    S => R1IN_ADD_1_1_AXB_10,
    LO => R1IN_ADD_1_1_CRY_10);
R1IN_ADD_1_1_S_9: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_9,
    CI => R1IN_ADD_1_1_CRY_8,
    O => N_1555);
R1IN_ADD_1_1_CRY_9_Z8017: MUXCY_L port map (
    DI => R1IN_3(41),
    CI => R1IN_ADD_1_1_CRY_8,
    S => R1IN_ADD_1_1_AXB_9,
    LO => R1IN_ADD_1_1_CRY_9);
R1IN_ADD_1_1_S_8: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_8,
    CI => R1IN_ADD_1_1_CRY_7,
    O => N_1553);
R1IN_ADD_1_1_CRY_8_Z8019: MUXCY_L port map (
    DI => R1IN_3(40),
    CI => R1IN_ADD_1_1_CRY_7,
    S => R1IN_ADD_1_1_AXB_8,
    LO => R1IN_ADD_1_1_CRY_8);
R1IN_ADD_1_1_S_7: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_7,
    CI => R1IN_ADD_1_1_CRY_6,
    O => N_1551);
R1IN_ADD_1_1_CRY_7_Z8021: MUXCY_L port map (
    DI => R1IN_3(39),
    CI => R1IN_ADD_1_1_CRY_6,
    S => R1IN_ADD_1_1_AXB_7,
    LO => R1IN_ADD_1_1_CRY_7);
R1IN_ADD_1_1_S_6: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_6,
    CI => R1IN_ADD_1_1_CRY_5,
    O => N_1549);
R1IN_ADD_1_1_CRY_6_Z8023: MUXCY_L port map (
    DI => R1IN_3(38),
    CI => R1IN_ADD_1_1_CRY_5,
    S => R1IN_ADD_1_1_AXB_6,
    LO => R1IN_ADD_1_1_CRY_6);
R1IN_ADD_1_1_S_5: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_5,
    CI => R1IN_ADD_1_1_CRY_4,
    O => N_1547);
R1IN_ADD_1_1_CRY_5_Z8025: MUXCY_L port map (
    DI => R1IN_3(37),
    CI => R1IN_ADD_1_1_CRY_4,
    S => R1IN_ADD_1_1_AXB_5,
    LO => R1IN_ADD_1_1_CRY_5);
R1IN_ADD_1_1_S_4: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_4,
    CI => R1IN_ADD_1_1_CRY_3,
    O => N_1545);
R1IN_ADD_1_1_CRY_4_Z8027: MUXCY_L port map (
    DI => R1IN_3(36),
    CI => R1IN_ADD_1_1_CRY_3,
    S => R1IN_ADD_1_1_AXB_4,
    LO => R1IN_ADD_1_1_CRY_4);
R1IN_ADD_1_1_S_3: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_3,
    CI => R1IN_ADD_1_1_CRY_2,
    O => N_1543);
R1IN_ADD_1_1_CRY_3_Z8029: MUXCY_L port map (
    DI => R1IN_3(35),
    CI => R1IN_ADD_1_1_CRY_2,
    S => R1IN_ADD_1_1_AXB_3,
    LO => R1IN_ADD_1_1_CRY_3);
R1IN_ADD_1_1_S_2: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_2,
    CI => R1IN_ADD_1_1_CRY_1,
    O => N_1541);
R1IN_ADD_1_1_CRY_2_Z8031: MUXCY_L port map (
    DI => R1IN_3(34),
    CI => R1IN_ADD_1_1_CRY_1,
    S => R1IN_ADD_1_1_AXB_2,
    LO => R1IN_ADD_1_1_CRY_2);
R1IN_ADD_1_1_S_1: XORCY port map (
    LI => R1IN_ADD_1_1_AXB_1,
    CI => R1IN_ADD_1_1_CRY_0,
    O => N_1539);
R1IN_ADD_1_1_CRY_1_Z8033: MUXCY_L port map (
    DI => R1IN_3(33),
    CI => R1IN_ADD_1_1_CRY_0,
    S => R1IN_ADD_1_1_AXB_1,
    LO => R1IN_ADD_1_1_CRY_1);
R1IN_ADD_1_1_CRY_0_Z8034: MUXCY_L port map (
    DI => R1IN_3(32),
    CI => NN_1,
    S => R1IN_ADD_1_1_AXB_0,
    LO => R1IN_ADD_1_1_CRY_0);
R1IN_ADD_1_0_S_31: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_31,
    CI => R1IN_ADD_1_0_CRY_30,
    O => R1IN_ADD_1(31));
R1IN_ADD_1_0_CRY_31_Z8036: MUXCY port map (
    DI => R1IN_3(31),
    CI => R1IN_ADD_1_0_CRY_30,
    S => R1IN_ADD_1_0_AXB_31,
    O => R1IN_ADD_1_0_CRY_31);
R1IN_ADD_1_0_S_30: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_30,
    CI => R1IN_ADD_1_0_CRY_29,
    O => R1IN_ADD_1(30));
R1IN_ADD_1_0_CRY_30_Z8038: MUXCY_L port map (
    DI => R1IN_3(30),
    CI => R1IN_ADD_1_0_CRY_29,
    S => R1IN_ADD_1_0_AXB_30,
    LO => R1IN_ADD_1_0_CRY_30);
R1IN_ADD_1_0_S_29: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_29,
    CI => R1IN_ADD_1_0_CRY_28,
    O => R1IN_ADD_1(29));
R1IN_ADD_1_0_CRY_29_Z8040: MUXCY_L port map (
    DI => R1IN_3(29),
    CI => R1IN_ADD_1_0_CRY_28,
    S => R1IN_ADD_1_0_AXB_29,
    LO => R1IN_ADD_1_0_CRY_29);
R1IN_ADD_1_0_S_28: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_28,
    CI => R1IN_ADD_1_0_CRY_27,
    O => R1IN_ADD_1(28));
R1IN_ADD_1_0_CRY_28_Z8042: MUXCY_L port map (
    DI => R1IN_3(28),
    CI => R1IN_ADD_1_0_CRY_27,
    S => R1IN_ADD_1_0_AXB_28,
    LO => R1IN_ADD_1_0_CRY_28);
R1IN_ADD_1_0_S_27: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_27,
    CI => R1IN_ADD_1_0_CRY_26,
    O => R1IN_ADD_1(27));
R1IN_ADD_1_0_CRY_27_Z8044: MUXCY_L port map (
    DI => R1IN_3(27),
    CI => R1IN_ADD_1_0_CRY_26,
    S => R1IN_ADD_1_0_AXB_27,
    LO => R1IN_ADD_1_0_CRY_27);
R1IN_ADD_1_0_S_26: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_26,
    CI => R1IN_ADD_1_0_CRY_25,
    O => R1IN_ADD_1(26));
R1IN_ADD_1_0_CRY_26_Z8046: MUXCY_L port map (
    DI => R1IN_3(26),
    CI => R1IN_ADD_1_0_CRY_25,
    S => R1IN_ADD_1_0_AXB_26,
    LO => R1IN_ADD_1_0_CRY_26);
R1IN_ADD_1_0_S_25: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_25,
    CI => R1IN_ADD_1_0_CRY_24,
    O => R1IN_ADD_1(25));
R1IN_ADD_1_0_CRY_25_Z8048: MUXCY_L port map (
    DI => R1IN_3(25),
    CI => R1IN_ADD_1_0_CRY_24,
    S => R1IN_ADD_1_0_AXB_25,
    LO => R1IN_ADD_1_0_CRY_25);
R1IN_ADD_1_0_S_24: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_24,
    CI => R1IN_ADD_1_0_CRY_23,
    O => R1IN_ADD_1(24));
R1IN_ADD_1_0_CRY_24_Z8050: MUXCY_L port map (
    DI => R1IN_3(24),
    CI => R1IN_ADD_1_0_CRY_23,
    S => R1IN_ADD_1_0_AXB_24,
    LO => R1IN_ADD_1_0_CRY_24);
R1IN_ADD_1_0_S_23: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_23,
    CI => R1IN_ADD_1_0_CRY_22,
    O => R1IN_ADD_1(23));
R1IN_ADD_1_0_CRY_23_Z8052: MUXCY_L port map (
    DI => R1IN_3(23),
    CI => R1IN_ADD_1_0_CRY_22,
    S => R1IN_ADD_1_0_AXB_23,
    LO => R1IN_ADD_1_0_CRY_23);
R1IN_ADD_1_0_S_22: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_22,
    CI => R1IN_ADD_1_0_CRY_21,
    O => R1IN_ADD_1(22));
R1IN_ADD_1_0_CRY_22_Z8054: MUXCY_L port map (
    DI => R1IN_3(22),
    CI => R1IN_ADD_1_0_CRY_21,
    S => R1IN_ADD_1_0_AXB_22,
    LO => R1IN_ADD_1_0_CRY_22);
R1IN_ADD_1_0_S_21: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_21,
    CI => R1IN_ADD_1_0_CRY_20,
    O => R1IN_ADD_1(21));
R1IN_ADD_1_0_CRY_21_Z8056: MUXCY_L port map (
    DI => R1IN_3(21),
    CI => R1IN_ADD_1_0_CRY_20,
    S => R1IN_ADD_1_0_AXB_21,
    LO => R1IN_ADD_1_0_CRY_21);
R1IN_ADD_1_0_S_20: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_20,
    CI => R1IN_ADD_1_0_CRY_19,
    O => R1IN_ADD_1(20));
R1IN_ADD_1_0_CRY_20_Z8058: MUXCY_L port map (
    DI => R1IN_3(20),
    CI => R1IN_ADD_1_0_CRY_19,
    S => R1IN_ADD_1_0_AXB_20,
    LO => R1IN_ADD_1_0_CRY_20);
R1IN_ADD_1_0_S_19: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_19,
    CI => R1IN_ADD_1_0_CRY_18,
    O => R1IN_ADD_1(19));
R1IN_ADD_1_0_CRY_19_Z8060: MUXCY_L port map (
    DI => R1IN_3(19),
    CI => R1IN_ADD_1_0_CRY_18,
    S => R1IN_ADD_1_0_AXB_19,
    LO => R1IN_ADD_1_0_CRY_19);
R1IN_ADD_1_0_S_18: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_18,
    CI => R1IN_ADD_1_0_CRY_17,
    O => R1IN_ADD_1(18));
R1IN_ADD_1_0_CRY_18_Z8062: MUXCY_L port map (
    DI => R1IN_3(18),
    CI => R1IN_ADD_1_0_CRY_17,
    S => R1IN_ADD_1_0_AXB_18,
    LO => R1IN_ADD_1_0_CRY_18);
R1IN_ADD_1_0_S_17: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_17,
    CI => R1IN_ADD_1_0_CRY_16,
    O => R1IN_ADD_1(17));
R1IN_ADD_1_0_CRY_17_Z8064: MUXCY_L port map (
    DI => R1IN_3(17),
    CI => R1IN_ADD_1_0_CRY_16,
    S => R1IN_ADD_1_0_AXB_17,
    LO => R1IN_ADD_1_0_CRY_17);
R1IN_ADD_1_0_S_16: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_16,
    CI => R1IN_ADD_1_0_CRY_15,
    O => R1IN_ADD_1(16));
R1IN_ADD_1_0_CRY_16_Z8066: MUXCY_L port map (
    DI => R1IN_2F(16),
    CI => R1IN_ADD_1_0_CRY_15,
    S => R1IN_ADD_1_0_AXB_16,
    LO => R1IN_ADD_1_0_CRY_16);
R1IN_ADD_1_0_S_15: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_15,
    CI => R1IN_ADD_1_0_CRY_14,
    O => R1IN_ADD_1(15));
R1IN_ADD_1_0_CRY_15_Z8068: MUXCY_L port map (
    DI => R1IN_2F(15),
    CI => R1IN_ADD_1_0_CRY_14,
    S => R1IN_ADD_1_0_AXB_15,
    LO => R1IN_ADD_1_0_CRY_15);
R1IN_ADD_1_0_S_14: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_14,
    CI => R1IN_ADD_1_0_CRY_13,
    O => R1IN_ADD_1(14));
R1IN_ADD_1_0_CRY_14_Z8070: MUXCY_L port map (
    DI => R1IN_2F(14),
    CI => R1IN_ADD_1_0_CRY_13,
    S => R1IN_ADD_1_0_AXB_14,
    LO => R1IN_ADD_1_0_CRY_14);
R1IN_ADD_1_0_S_13: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_13,
    CI => R1IN_ADD_1_0_CRY_12,
    O => R1IN_ADD_1(13));
R1IN_ADD_1_0_CRY_13_Z8072: MUXCY_L port map (
    DI => R1IN_2F(13),
    CI => R1IN_ADD_1_0_CRY_12,
    S => R1IN_ADD_1_0_AXB_13,
    LO => R1IN_ADD_1_0_CRY_13);
R1IN_ADD_1_0_S_12: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_12,
    CI => R1IN_ADD_1_0_CRY_11,
    O => R1IN_ADD_1(12));
R1IN_ADD_1_0_CRY_12_Z8074: MUXCY_L port map (
    DI => R1IN_2F(12),
    CI => R1IN_ADD_1_0_CRY_11,
    S => R1IN_ADD_1_0_AXB_12,
    LO => R1IN_ADD_1_0_CRY_12);
R1IN_ADD_1_0_S_11: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_11,
    CI => R1IN_ADD_1_0_CRY_10,
    O => R1IN_ADD_1(11));
R1IN_ADD_1_0_CRY_11_Z8076: MUXCY_L port map (
    DI => R1IN_2F(11),
    CI => R1IN_ADD_1_0_CRY_10,
    S => R1IN_ADD_1_0_AXB_11,
    LO => R1IN_ADD_1_0_CRY_11);
R1IN_ADD_1_0_S_10: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_10,
    CI => R1IN_ADD_1_0_CRY_9,
    O => R1IN_ADD_1(10));
R1IN_ADD_1_0_CRY_10_Z8078: MUXCY_L port map (
    DI => R1IN_2F(10),
    CI => R1IN_ADD_1_0_CRY_9,
    S => R1IN_ADD_1_0_AXB_10,
    LO => R1IN_ADD_1_0_CRY_10);
R1IN_ADD_1_0_S_9: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_9,
    CI => R1IN_ADD_1_0_CRY_8,
    O => R1IN_ADD_1(9));
R1IN_ADD_1_0_CRY_9_Z8080: MUXCY_L port map (
    DI => R1IN_2F(9),
    CI => R1IN_ADD_1_0_CRY_8,
    S => R1IN_ADD_1_0_AXB_9,
    LO => R1IN_ADD_1_0_CRY_9);
R1IN_ADD_1_0_S_8: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_8,
    CI => R1IN_ADD_1_0_CRY_7,
    O => R1IN_ADD_1(8));
R1IN_ADD_1_0_CRY_8_Z8082: MUXCY_L port map (
    DI => R1IN_2F(8),
    CI => R1IN_ADD_1_0_CRY_7,
    S => R1IN_ADD_1_0_AXB_8,
    LO => R1IN_ADD_1_0_CRY_8);
R1IN_ADD_1_0_S_7: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_7,
    CI => R1IN_ADD_1_0_CRY_6,
    O => R1IN_ADD_1(7));
R1IN_ADD_1_0_CRY_7_Z8084: MUXCY_L port map (
    DI => R1IN_2F(7),
    CI => R1IN_ADD_1_0_CRY_6,
    S => R1IN_ADD_1_0_AXB_7,
    LO => R1IN_ADD_1_0_CRY_7);
R1IN_ADD_1_0_S_6: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_6,
    CI => R1IN_ADD_1_0_CRY_5,
    O => R1IN_ADD_1(6));
R1IN_ADD_1_0_CRY_6_Z8086: MUXCY_L port map (
    DI => R1IN_2F(6),
    CI => R1IN_ADD_1_0_CRY_5,
    S => R1IN_ADD_1_0_AXB_6,
    LO => R1IN_ADD_1_0_CRY_6);
R1IN_ADD_1_0_S_5: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_5,
    CI => R1IN_ADD_1_0_CRY_4,
    O => R1IN_ADD_1(5));
R1IN_ADD_1_0_CRY_5_Z8088: MUXCY_L port map (
    DI => R1IN_2F(5),
    CI => R1IN_ADD_1_0_CRY_4,
    S => R1IN_ADD_1_0_AXB_5,
    LO => R1IN_ADD_1_0_CRY_5);
R1IN_ADD_1_0_S_4: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_4,
    CI => R1IN_ADD_1_0_CRY_3,
    O => R1IN_ADD_1(4));
R1IN_ADD_1_0_CRY_4_Z8090: MUXCY_L port map (
    DI => R1IN_2F(4),
    CI => R1IN_ADD_1_0_CRY_3,
    S => R1IN_ADD_1_0_AXB_4,
    LO => R1IN_ADD_1_0_CRY_4);
R1IN_ADD_1_0_S_3: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_3,
    CI => R1IN_ADD_1_0_CRY_2,
    O => R1IN_ADD_1(3));
R1IN_ADD_1_0_CRY_3_Z8092: MUXCY_L port map (
    DI => R1IN_2F(3),
    CI => R1IN_ADD_1_0_CRY_2,
    S => R1IN_ADD_1_0_AXB_3,
    LO => R1IN_ADD_1_0_CRY_3);
R1IN_ADD_1_0_S_2: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_2,
    CI => R1IN_ADD_1_0_CRY_1,
    O => R1IN_ADD_1(2));
R1IN_ADD_1_0_CRY_2_Z8094: MUXCY_L port map (
    DI => R1IN_2F(2),
    CI => R1IN_ADD_1_0_CRY_1,
    S => R1IN_ADD_1_0_AXB_2,
    LO => R1IN_ADD_1_0_CRY_2);
R1IN_ADD_1_0_S_1: XORCY port map (
    LI => R1IN_ADD_1_0_AXB_1,
    CI => R1IN_ADD_1_0_CRY_0,
    O => R1IN_ADD_1(1));
R1IN_ADD_1_0_CRY_1_Z8096: MUXCY_L port map (
    DI => R1IN_2F(1),
    CI => R1IN_ADD_1_0_CRY_0,
    S => R1IN_ADD_1_0_AXB_1,
    LO => R1IN_ADD_1_0_CRY_1);
R1IN_ADD_1_0_CRY_0_Z8097: MUXCY_L port map (
    DI => R1IN_2F(0),
    CI => NN_1,
    S => R1IN_ADD_1(0),
    LO => R1IN_ADD_1_0_CRY_0);
R1IN_ADD_2_1_0_S_51_Z8098: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_51,
    CI => R1IN_ADD_2_1_0_CRY_50,
    O => R1IN_ADD_2_1_0_S_51);
R1IN_ADD_2_1_0_S_50_Z8099: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_50,
    CI => R1IN_ADD_2_1_0_CRY_49,
    O => R1IN_ADD_2_1_0_S_50);
R1IN_ADD_2_1_0_CRY_50_Z8100: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_49,
    S => R1IN_ADD_2_1_0_AXB_50,
    LO => R1IN_ADD_2_1_0_CRY_50);
R1IN_ADD_2_1_0_S_49_Z8101: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_49,
    CI => R1IN_ADD_2_1_0_CRY_48,
    O => R1IN_ADD_2_1_0_S_49);
R1IN_ADD_2_1_0_CRY_49_Z8102: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_48,
    S => R1IN_ADD_2_1_0_AXB_49,
    LO => R1IN_ADD_2_1_0_CRY_49);
R1IN_ADD_2_1_0_S_48_Z8103: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_48,
    CI => R1IN_ADD_2_1_0_CRY_47,
    O => R1IN_ADD_2_1_0_S_48);
R1IN_ADD_2_1_0_CRY_48_Z8104: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_47,
    S => R1IN_ADD_2_1_0_AXB_48,
    LO => R1IN_ADD_2_1_0_CRY_48);
R1IN_ADD_2_1_0_S_47_Z8105: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_47,
    CI => R1IN_ADD_2_1_0_CRY_46,
    O => R1IN_ADD_2_1_0_S_47);
R1IN_ADD_2_1_0_CRY_47_Z8106: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_46,
    S => R1IN_ADD_2_1_0_AXB_47,
    LO => R1IN_ADD_2_1_0_CRY_47);
R1IN_ADD_2_1_0_S_46_Z8107: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_46,
    CI => R1IN_ADD_2_1_0_CRY_45,
    O => R1IN_ADD_2_1_0_S_46);
R1IN_ADD_2_1_0_CRY_46_Z8108: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_45,
    S => R1IN_ADD_2_1_0_AXB_46,
    LO => R1IN_ADD_2_1_0_CRY_46);
R1IN_ADD_2_1_0_S_45_Z8109: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_45,
    CI => R1IN_ADD_2_1_0_CRY_44,
    O => R1IN_ADD_2_1_0_S_45);
R1IN_ADD_2_1_0_CRY_45_Z8110: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_44,
    S => R1IN_ADD_2_1_0_AXB_45,
    LO => R1IN_ADD_2_1_0_CRY_45);
R1IN_ADD_2_1_0_S_44_Z8111: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_44,
    CI => R1IN_ADD_2_1_0_CRY_43,
    O => R1IN_ADD_2_1_0_S_44);
R1IN_ADD_2_1_0_CRY_44_Z8112: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_43,
    S => R1IN_ADD_2_1_0_AXB_44,
    LO => R1IN_ADD_2_1_0_CRY_44);
R1IN_ADD_2_1_0_S_43_Z8113: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_43,
    CI => R1IN_ADD_2_1_0_CRY_42,
    O => R1IN_ADD_2_1_0_S_43);
R1IN_ADD_2_1_0_CRY_43_Z8114: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_42,
    S => R1IN_ADD_2_1_0_AXB_43,
    LO => R1IN_ADD_2_1_0_CRY_43);
R1IN_ADD_2_1_0_S_42_Z8115: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_42,
    CI => R1IN_ADD_2_1_0_CRY_41,
    O => R1IN_ADD_2_1_0_S_42);
R1IN_ADD_2_1_0_CRY_42_Z8116: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_41,
    S => R1IN_ADD_2_1_0_AXB_42,
    LO => R1IN_ADD_2_1_0_CRY_42);
R1IN_ADD_2_1_0_S_41_Z8117: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_41,
    CI => R1IN_ADD_2_1_0_CRY_40,
    O => R1IN_ADD_2_1_0_S_41);
R1IN_ADD_2_1_0_CRY_41_Z8118: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_40,
    S => R1IN_ADD_2_1_0_AXB_41,
    LO => R1IN_ADD_2_1_0_CRY_41);
R1IN_ADD_2_1_0_S_40_Z8119: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_40,
    CI => R1IN_ADD_2_1_0_CRY_39,
    O => R1IN_ADD_2_1_0_S_40);
R1IN_ADD_2_1_0_CRY_40_Z8120: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_39,
    S => R1IN_ADD_2_1_0_AXB_40,
    LO => R1IN_ADD_2_1_0_CRY_40);
R1IN_ADD_2_1_0_S_39_Z8121: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_39,
    CI => R1IN_ADD_2_1_0_CRY_38,
    O => R1IN_ADD_2_1_0_S_39);
R1IN_ADD_2_1_0_CRY_39_Z8122: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_38,
    S => R1IN_ADD_2_1_0_AXB_39,
    LO => R1IN_ADD_2_1_0_CRY_39);
R1IN_ADD_2_1_0_S_38_Z8123: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_38,
    CI => R1IN_ADD_2_1_0_CRY_37,
    O => R1IN_ADD_2_1_0_S_38);
R1IN_ADD_2_1_0_CRY_38_Z8124: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_37,
    S => R1IN_ADD_2_1_0_AXB_38,
    LO => R1IN_ADD_2_1_0_CRY_38);
R1IN_ADD_2_1_0_S_37_Z8125: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_37,
    CI => R1IN_ADD_2_1_0_CRY_36,
    O => R1IN_ADD_2_1_0_S_37);
R1IN_ADD_2_1_0_CRY_37_Z8126: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_36,
    S => R1IN_ADD_2_1_0_AXB_37,
    LO => R1IN_ADD_2_1_0_CRY_37);
R1IN_ADD_2_1_0_S_36_Z8127: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_36,
    CI => R1IN_ADD_2_1_0_CRY_35,
    O => R1IN_ADD_2_1_0_S_36);
R1IN_ADD_2_1_0_CRY_36_Z8128: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_35,
    S => R1IN_ADD_2_1_0_AXB_36,
    LO => R1IN_ADD_2_1_0_CRY_36);
R1IN_ADD_2_1_0_S_35_Z8129: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_35,
    CI => R1IN_ADD_2_1_0_CRY_34,
    O => R1IN_ADD_2_1_0_S_35);
R1IN_ADD_2_1_0_CRY_35_Z8130: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_34,
    S => R1IN_ADD_2_1_0_AXB_35,
    LO => R1IN_ADD_2_1_0_CRY_35);
R1IN_ADD_2_1_0_S_34_Z8131: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_34,
    CI => R1IN_ADD_2_1_0_CRY_33,
    O => R1IN_ADD_2_1_0_S_34);
R1IN_ADD_2_1_0_CRY_34_Z8132: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_33,
    S => R1IN_ADD_2_1_0_AXB_34,
    LO => R1IN_ADD_2_1_0_CRY_34);
R1IN_ADD_2_1_0_S_33_Z8133: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_33,
    CI => R1IN_ADD_2_1_0_CRY_32,
    O => R1IN_ADD_2_1_0_S_33);
R1IN_ADD_2_1_0_CRY_33_Z8134: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_32,
    S => R1IN_ADD_2_1_0_AXB_33,
    LO => R1IN_ADD_2_1_0_CRY_33);
R1IN_ADD_2_1_0_S_32_Z8135: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_32,
    CI => R1IN_ADD_2_1_0_CRY_31,
    O => R1IN_ADD_2_1_0_S_32);
R1IN_ADD_2_1_0_CRY_32_Z8136: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_31,
    S => R1IN_ADD_2_1_0_AXB_32,
    LO => R1IN_ADD_2_1_0_CRY_32);
R1IN_ADD_2_1_0_S_31_Z8137: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_31,
    CI => R1IN_ADD_2_1_0_CRY_30,
    O => R1IN_ADD_2_1_0_S_31);
R1IN_ADD_2_1_0_CRY_31_Z8138: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_30,
    S => R1IN_ADD_2_1_0_AXB_31,
    LO => R1IN_ADD_2_1_0_CRY_31);
R1IN_ADD_2_1_0_S_30_Z8139: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_30,
    CI => R1IN_ADD_2_1_0_CRY_29,
    O => R1IN_ADD_2_1_0_S_30);
R1IN_ADD_2_1_0_CRY_30_Z8140: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_29,
    S => R1IN_ADD_2_1_0_AXB_30,
    LO => R1IN_ADD_2_1_0_CRY_30);
R1IN_ADD_2_1_0_S_29_Z8141: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_29,
    CI => R1IN_ADD_2_1_0_CRY_28,
    O => R1IN_ADD_2_1_0_S_29);
R1IN_ADD_2_1_0_CRY_29_Z8142: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_28,
    S => R1IN_ADD_2_1_0_AXB_29,
    LO => R1IN_ADD_2_1_0_CRY_29);
R1IN_ADD_2_1_0_S_28_Z8143: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_28,
    CI => R1IN_ADD_2_1_0_CRY_27,
    O => R1IN_ADD_2_1_0_S_28);
R1IN_ADD_2_1_0_CRY_28_Z8144: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_27,
    S => R1IN_ADD_2_1_0_AXB_28,
    LO => R1IN_ADD_2_1_0_CRY_28);
R1IN_ADD_2_1_0_S_27_Z8145: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_27,
    CI => R1IN_ADD_2_1_0_CRY_26,
    O => R1IN_ADD_2_1_0_S_27);
R1IN_ADD_2_1_0_CRY_27_Z8146: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_26,
    S => R1IN_ADD_2_1_0_AXB_27,
    LO => R1IN_ADD_2_1_0_CRY_27);
R1IN_ADD_2_1_0_S_26_Z8147: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_26,
    CI => R1IN_ADD_2_1_0_CRY_25,
    O => R1IN_ADD_2_1_0_S_26);
R1IN_ADD_2_1_0_CRY_26_Z8148: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_25,
    S => R1IN_ADD_2_1_0_AXB_26,
    LO => R1IN_ADD_2_1_0_CRY_26);
R1IN_ADD_2_1_0_S_25_Z8149: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_25,
    CI => R1IN_ADD_2_1_0_CRY_24,
    O => R1IN_ADD_2_1_0_S_25);
R1IN_ADD_2_1_0_CRY_25_Z8150: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_24,
    S => R1IN_ADD_2_1_0_AXB_25,
    LO => R1IN_ADD_2_1_0_CRY_25);
R1IN_ADD_2_1_0_S_24_Z8151: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_24,
    CI => R1IN_ADD_2_1_0_CRY_23,
    O => R1IN_ADD_2_1_0_S_24);
R1IN_ADD_2_1_0_CRY_24_Z8152: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_23,
    S => R1IN_ADD_2_1_0_AXB_24,
    LO => R1IN_ADD_2_1_0_CRY_24);
R1IN_ADD_2_1_0_S_23_Z8153: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_23,
    CI => R1IN_ADD_2_1_0_CRY_22,
    O => R1IN_ADD_2_1_0_S_23);
R1IN_ADD_2_1_0_CRY_23_Z8154: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_22,
    S => R1IN_ADD_2_1_0_AXB_23,
    LO => R1IN_ADD_2_1_0_CRY_23);
R1IN_ADD_2_1_0_S_22_Z8155: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_22,
    CI => R1IN_ADD_2_1_0_CRY_21,
    O => R1IN_ADD_2_1_0_S_22);
R1IN_ADD_2_1_0_CRY_22_Z8156: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_21,
    S => R1IN_ADD_2_1_0_AXB_22,
    LO => R1IN_ADD_2_1_0_CRY_22);
R1IN_ADD_2_1_0_S_21_Z8157: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_21,
    CI => R1IN_ADD_2_1_0_CRY_20,
    O => R1IN_ADD_2_1_0_S_21);
R1IN_ADD_2_1_0_CRY_21_Z8158: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_20,
    S => R1IN_ADD_2_1_0_AXB_21,
    LO => R1IN_ADD_2_1_0_CRY_21);
R1IN_ADD_2_1_0_S_20_Z8159: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_20,
    CI => R1IN_ADD_2_1_0_CRY_19,
    O => R1IN_ADD_2_1_0_S_20);
R1IN_ADD_2_1_0_CRY_20_Z8160: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_19,
    S => R1IN_ADD_2_1_0_AXB_20,
    LO => R1IN_ADD_2_1_0_CRY_20);
R1IN_ADD_2_1_0_S_19_Z8161: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_19,
    CI => R1IN_ADD_2_1_0_CRY_18,
    O => R1IN_ADD_2_1_0_S_19);
R1IN_ADD_2_1_0_CRY_19_Z8162: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_18,
    S => R1IN_ADD_2_1_0_AXB_19,
    LO => R1IN_ADD_2_1_0_CRY_19);
R1IN_ADD_2_1_0_S_18_Z8163: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_18,
    CI => R1IN_ADD_2_1_0_CRY_17,
    O => R1IN_ADD_2_1_0_S_18);
R1IN_ADD_2_1_0_CRY_18_Z8164: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_17,
    S => R1IN_ADD_2_1_0_AXB_18,
    LO => R1IN_ADD_2_1_0_CRY_18);
R1IN_ADD_2_1_0_S_17_Z8165: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_17,
    CI => R1IN_ADD_2_1_0_CRY_16,
    O => R1IN_ADD_2_1_0_S_17);
R1IN_ADD_2_1_0_CRY_17_Z8166: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_16,
    S => R1IN_ADD_2_1_0_AXB_17,
    LO => R1IN_ADD_2_1_0_CRY_17);
R1IN_ADD_2_1_0_S_16_Z8167: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_16,
    CI => R1IN_ADD_2_1_0_CRY_15,
    O => R1IN_ADD_2_1_0_S_16);
R1IN_ADD_2_1_0_CRY_16_Z8168: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_15,
    S => R1IN_ADD_2_1_0_AXB_16,
    LO => R1IN_ADD_2_1_0_CRY_16);
R1IN_ADD_2_1_0_S_15_Z8169: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_15,
    CI => R1IN_ADD_2_1_0_CRY_14,
    O => R1IN_ADD_2_1_0_S_15);
R1IN_ADD_2_1_0_CRY_15_Z8170: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_14,
    S => R1IN_ADD_2_1_0_AXB_15,
    LO => R1IN_ADD_2_1_0_CRY_15);
R1IN_ADD_2_1_0_S_14_Z8171: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_14,
    CI => R1IN_ADD_2_1_0_CRY_13,
    O => R1IN_ADD_2_1_0_S_14);
R1IN_ADD_2_1_0_CRY_14_Z8172: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_13,
    S => R1IN_ADD_2_1_0_AXB_14,
    LO => R1IN_ADD_2_1_0_CRY_14);
R1IN_ADD_2_1_0_S_13_Z8173: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_13,
    CI => R1IN_ADD_2_1_0_CRY_12,
    O => R1IN_ADD_2_1_0_S_13);
R1IN_ADD_2_1_0_CRY_13_Z8174: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_12,
    S => R1IN_ADD_2_1_0_AXB_13,
    LO => R1IN_ADD_2_1_0_CRY_13);
R1IN_ADD_2_1_0_S_12_Z8175: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_12,
    CI => R1IN_ADD_2_1_0_CRY_11,
    O => R1IN_ADD_2_1_0_S_12);
R1IN_ADD_2_1_0_CRY_12_Z8176: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_11,
    S => R1IN_ADD_2_1_0_AXB_12,
    LO => R1IN_ADD_2_1_0_CRY_12);
R1IN_ADD_2_1_0_S_11_Z8177: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_11,
    CI => R1IN_ADD_2_1_0_CRY_10,
    O => R1IN_ADD_2_1_0_S_11);
R1IN_ADD_2_1_0_CRY_11_Z8178: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_10,
    S => R1IN_ADD_2_1_0_AXB_11,
    LO => R1IN_ADD_2_1_0_CRY_11);
R1IN_ADD_2_1_0_S_10_Z8179: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_10,
    CI => R1IN_ADD_2_1_0_CRY_9,
    O => R1IN_ADD_2_1_0_S_10);
R1IN_ADD_2_1_0_CRY_10_Z8180: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_9,
    S => R1IN_ADD_2_1_0_AXB_10,
    LO => R1IN_ADD_2_1_0_CRY_10);
R1IN_ADD_2_1_0_S_9_Z8181: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_9,
    CI => R1IN_ADD_2_1_0_CRY_8,
    O => R1IN_ADD_2_1_0_S_9);
R1IN_ADD_2_1_0_CRY_9_Z8182: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_0_CRY_8,
    S => R1IN_ADD_2_1_0_AXB_9,
    LO => R1IN_ADD_2_1_0_CRY_9);
R1IN_ADD_2_1_0_S_8_Z8183: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_8,
    CI => R1IN_ADD_2_1_0_CRY_7,
    O => R1IN_ADD_2_1_0_S_8);
R1IN_ADD_2_1_0_CRY_8_Z8184: MUXCY_L port map (
    DI => R1IN_4F(44),
    CI => R1IN_ADD_2_1_0_CRY_7,
    S => R1IN_ADD_2_1_0_AXB_8,
    LO => R1IN_ADD_2_1_0_CRY_8);
R1IN_ADD_2_1_0_S_7_Z8185: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_7,
    CI => R1IN_ADD_2_1_0_CRY_6,
    O => R1IN_ADD_2_1_0_S_7);
R1IN_ADD_2_1_0_CRY_7_Z8186: MUXCY_L port map (
    DI => R1IN_4F(43),
    CI => R1IN_ADD_2_1_0_CRY_6,
    S => R1IN_ADD_2_1_0_AXB_7,
    LO => R1IN_ADD_2_1_0_CRY_7);
R1IN_ADD_2_1_0_S_6_Z8187: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_6,
    CI => R1IN_ADD_2_1_0_CRY_5,
    O => R1IN_ADD_2_1_0_S_6);
R1IN_ADD_2_1_0_CRY_6_Z8188: MUXCY_L port map (
    DI => R1IN_4F(42),
    CI => R1IN_ADD_2_1_0_CRY_5,
    S => R1IN_ADD_2_1_0_AXB_6,
    LO => R1IN_ADD_2_1_0_CRY_6);
R1IN_ADD_2_1_0_S_5_Z8189: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_5,
    CI => R1IN_ADD_2_1_0_CRY_4,
    O => R1IN_ADD_2_1_0_S_5);
R1IN_ADD_2_1_0_CRY_5_Z8190: MUXCY_L port map (
    DI => R1IN_4F(41),
    CI => R1IN_ADD_2_1_0_CRY_4,
    S => R1IN_ADD_2_1_0_AXB_5,
    LO => R1IN_ADD_2_1_0_CRY_5);
R1IN_ADD_2_1_0_S_4_Z8191: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_4,
    CI => R1IN_ADD_2_1_0_CRY_3,
    O => R1IN_ADD_2_1_0_S_4);
R1IN_ADD_2_1_0_CRY_4_Z8192: MUXCY_L port map (
    DI => R1IN_4F(40),
    CI => R1IN_ADD_2_1_0_CRY_3,
    S => R1IN_ADD_2_1_0_AXB_4,
    LO => R1IN_ADD_2_1_0_CRY_4);
R1IN_ADD_2_1_0_S_3_Z8193: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_3,
    CI => R1IN_ADD_2_1_0_CRY_2,
    O => R1IN_ADD_2_1_0_S_3);
R1IN_ADD_2_1_0_CRY_3_Z8194: MUXCY_L port map (
    DI => R1IN_4F(39),
    CI => R1IN_ADD_2_1_0_CRY_2,
    S => R1IN_ADD_2_1_0_AXB_3,
    LO => R1IN_ADD_2_1_0_CRY_3);
R1IN_ADD_2_1_0_S_2_Z8195: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_2,
    CI => R1IN_ADD_2_1_0_CRY_1,
    O => R1IN_ADD_2_1_0_S_2);
R1IN_ADD_2_1_0_CRY_2_Z8196: MUXCY_L port map (
    DI => R1IN_4F(38),
    CI => R1IN_ADD_2_1_0_CRY_1,
    S => R1IN_ADD_2_1_0_AXB_2,
    LO => R1IN_ADD_2_1_0_CRY_2);
R1IN_ADD_2_1_0_S_1_Z8197: XORCY port map (
    LI => R1IN_ADD_2_1_0_AXB_1,
    CI => R1IN_ADD_2_1_0_CRY_0,
    O => R1IN_ADD_2_1_0_S_1);
R1IN_ADD_2_1_0_CRY_1_Z8198: MUXCY_L port map (
    DI => R1IN_4F(37),
    CI => R1IN_ADD_2_1_0_CRY_0,
    S => R1IN_ADD_2_1_0_AXB_1,
    LO => R1IN_ADD_2_1_0_CRY_1);
R1IN_ADD_2_1_0_CRY_0_Z8199: MUXCY_L port map (
    DI => R1IN_4F(36),
    CI => NN_2,
    S => R1IN_ADD_2_1_0_AXB_0,
    LO => R1IN_ADD_2_1_0_CRY_0);
R1IN_ADD_2_1_S_51_Z8200: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_51,
    CI => R1IN_ADD_2_1_CRY_50,
    O => R1IN_ADD_2_1_S_51);
R1IN_ADD_2_1_S_50_Z8201: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_50,
    CI => R1IN_ADD_2_1_CRY_49,
    O => R1IN_ADD_2_1_S_50);
R1IN_ADD_2_1_CRY_50_Z8202: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_49,
    S => R1IN_ADD_2_1_AXB_50,
    LO => R1IN_ADD_2_1_CRY_50);
R1IN_ADD_2_1_S_49_Z8203: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_49,
    CI => R1IN_ADD_2_1_CRY_48,
    O => R1IN_ADD_2_1_S_49);
R1IN_ADD_2_1_CRY_49_Z8204: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_48,
    S => R1IN_ADD_2_1_AXB_49,
    LO => R1IN_ADD_2_1_CRY_49);
R1IN_ADD_2_1_S_48_Z8205: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_48,
    CI => R1IN_ADD_2_1_CRY_47,
    O => R1IN_ADD_2_1_S_48);
R1IN_ADD_2_1_CRY_48_Z8206: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_47,
    S => R1IN_ADD_2_1_AXB_48,
    LO => R1IN_ADD_2_1_CRY_48);
R1IN_ADD_2_1_S_47_Z8207: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_47,
    CI => R1IN_ADD_2_1_CRY_46,
    O => R1IN_ADD_2_1_S_47);
R1IN_ADD_2_1_CRY_47_Z8208: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_46,
    S => R1IN_ADD_2_1_AXB_47,
    LO => R1IN_ADD_2_1_CRY_47);
R1IN_ADD_2_1_S_46_Z8209: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_46,
    CI => R1IN_ADD_2_1_CRY_45,
    O => R1IN_ADD_2_1_S_46);
R1IN_ADD_2_1_CRY_46_Z8210: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_45,
    S => R1IN_ADD_2_1_AXB_46,
    LO => R1IN_ADD_2_1_CRY_46);
R1IN_ADD_2_1_S_45_Z8211: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_45,
    CI => R1IN_ADD_2_1_CRY_44,
    O => R1IN_ADD_2_1_S_45);
R1IN_ADD_2_1_CRY_45_Z8212: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_44,
    S => R1IN_ADD_2_1_AXB_45,
    LO => R1IN_ADD_2_1_CRY_45);
R1IN_ADD_2_1_S_44_Z8213: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_44,
    CI => R1IN_ADD_2_1_CRY_43,
    O => R1IN_ADD_2_1_S_44);
R1IN_ADD_2_1_CRY_44_Z8214: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_43,
    S => R1IN_ADD_2_1_AXB_44,
    LO => R1IN_ADD_2_1_CRY_44);
R1IN_ADD_2_1_S_43_Z8215: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_43,
    CI => R1IN_ADD_2_1_CRY_42,
    O => R1IN_ADD_2_1_S_43);
R1IN_ADD_2_1_CRY_43_Z8216: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_42,
    S => R1IN_ADD_2_1_AXB_43,
    LO => R1IN_ADD_2_1_CRY_43);
R1IN_ADD_2_1_S_42_Z8217: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_42,
    CI => R1IN_ADD_2_1_CRY_41,
    O => R1IN_ADD_2_1_S_42);
R1IN_ADD_2_1_CRY_42_Z8218: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_41,
    S => R1IN_ADD_2_1_AXB_42,
    LO => R1IN_ADD_2_1_CRY_42);
R1IN_ADD_2_1_S_41_Z8219: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_41,
    CI => R1IN_ADD_2_1_CRY_40,
    O => R1IN_ADD_2_1_S_41);
R1IN_ADD_2_1_CRY_41_Z8220: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_40,
    S => R1IN_ADD_2_1_AXB_41,
    LO => R1IN_ADD_2_1_CRY_41);
R1IN_ADD_2_1_S_40_Z8221: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_40,
    CI => R1IN_ADD_2_1_CRY_39,
    O => R1IN_ADD_2_1_S_40);
R1IN_ADD_2_1_CRY_40_Z8222: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_39,
    S => R1IN_ADD_2_1_AXB_40,
    LO => R1IN_ADD_2_1_CRY_40);
R1IN_ADD_2_1_S_39_Z8223: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_39,
    CI => R1IN_ADD_2_1_CRY_38,
    O => R1IN_ADD_2_1_S_39);
R1IN_ADD_2_1_CRY_39_Z8224: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_38,
    S => R1IN_ADD_2_1_AXB_39,
    LO => R1IN_ADD_2_1_CRY_39);
R1IN_ADD_2_1_S_38_Z8225: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_38,
    CI => R1IN_ADD_2_1_CRY_37,
    O => R1IN_ADD_2_1_S_38);
R1IN_ADD_2_1_CRY_38_Z8226: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_37,
    S => R1IN_ADD_2_1_AXB_38,
    LO => R1IN_ADD_2_1_CRY_38);
R1IN_ADD_2_1_S_37_Z8227: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_37,
    CI => R1IN_ADD_2_1_CRY_36,
    O => R1IN_ADD_2_1_S_37);
R1IN_ADD_2_1_CRY_37_Z8228: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_36,
    S => R1IN_ADD_2_1_AXB_37,
    LO => R1IN_ADD_2_1_CRY_37);
R1IN_ADD_2_1_S_36_Z8229: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_36,
    CI => R1IN_ADD_2_1_CRY_35,
    O => R1IN_ADD_2_1_S_36);
R1IN_ADD_2_1_CRY_36_Z8230: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_35,
    S => R1IN_ADD_2_1_AXB_36,
    LO => R1IN_ADD_2_1_CRY_36);
R1IN_ADD_2_1_S_35_Z8231: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_35,
    CI => R1IN_ADD_2_1_CRY_34,
    O => R1IN_ADD_2_1_S_35);
R1IN_ADD_2_1_CRY_35_Z8232: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_34,
    S => R1IN_ADD_2_1_AXB_35,
    LO => R1IN_ADD_2_1_CRY_35);
R1IN_ADD_2_1_S_34_Z8233: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_34,
    CI => R1IN_ADD_2_1_CRY_33,
    O => R1IN_ADD_2_1_S_34);
R1IN_ADD_2_1_CRY_34_Z8234: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_33,
    S => R1IN_ADD_2_1_AXB_34,
    LO => R1IN_ADD_2_1_CRY_34);
R1IN_ADD_2_1_S_33_Z8235: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_33,
    CI => R1IN_ADD_2_1_CRY_32,
    O => R1IN_ADD_2_1_S_33);
R1IN_ADD_2_1_CRY_33_Z8236: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_32,
    S => R1IN_ADD_2_1_AXB_33,
    LO => R1IN_ADD_2_1_CRY_33);
R1IN_ADD_2_1_S_32_Z8237: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_32,
    CI => R1IN_ADD_2_1_CRY_31,
    O => R1IN_ADD_2_1_S_32);
R1IN_ADD_2_1_CRY_32_Z8238: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_31,
    S => R1IN_ADD_2_1_AXB_32,
    LO => R1IN_ADD_2_1_CRY_32);
R1IN_ADD_2_1_S_31_Z8239: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_31,
    CI => R1IN_ADD_2_1_CRY_30,
    O => R1IN_ADD_2_1_S_31);
R1IN_ADD_2_1_CRY_31_Z8240: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_30,
    S => R1IN_ADD_2_1_AXB_31,
    LO => R1IN_ADD_2_1_CRY_31);
R1IN_ADD_2_1_S_30_Z8241: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_30,
    CI => R1IN_ADD_2_1_CRY_29,
    O => R1IN_ADD_2_1_S_30);
R1IN_ADD_2_1_CRY_30_Z8242: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_29,
    S => R1IN_ADD_2_1_AXB_30,
    LO => R1IN_ADD_2_1_CRY_30);
R1IN_ADD_2_1_S_29_Z8243: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_29,
    CI => R1IN_ADD_2_1_CRY_28,
    O => R1IN_ADD_2_1_S_29);
R1IN_ADD_2_1_CRY_29_Z8244: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_28,
    S => R1IN_ADD_2_1_AXB_29,
    LO => R1IN_ADD_2_1_CRY_29);
R1IN_ADD_2_1_S_28_Z8245: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_28,
    CI => R1IN_ADD_2_1_CRY_27,
    O => R1IN_ADD_2_1_S_28);
R1IN_ADD_2_1_CRY_28_Z8246: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_27,
    S => R1IN_ADD_2_1_AXB_28,
    LO => R1IN_ADD_2_1_CRY_28);
R1IN_ADD_2_1_S_27_Z8247: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_27,
    CI => R1IN_ADD_2_1_CRY_26,
    O => R1IN_ADD_2_1_S_27);
R1IN_ADD_2_1_CRY_27_Z8248: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_26,
    S => R1IN_ADD_2_1_AXB_27,
    LO => R1IN_ADD_2_1_CRY_27);
R1IN_ADD_2_1_S_26_Z8249: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_26,
    CI => R1IN_ADD_2_1_CRY_25,
    O => R1IN_ADD_2_1_S_26);
R1IN_ADD_2_1_CRY_26_Z8250: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_25,
    S => R1IN_ADD_2_1_AXB_26,
    LO => R1IN_ADD_2_1_CRY_26);
R1IN_ADD_2_1_S_25_Z8251: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_25,
    CI => R1IN_ADD_2_1_CRY_24,
    O => R1IN_ADD_2_1_S_25);
R1IN_ADD_2_1_CRY_25_Z8252: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_24,
    S => R1IN_ADD_2_1_AXB_25,
    LO => R1IN_ADD_2_1_CRY_25);
R1IN_ADD_2_1_S_24_Z8253: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_24,
    CI => R1IN_ADD_2_1_CRY_23,
    O => R1IN_ADD_2_1_S_24);
R1IN_ADD_2_1_CRY_24_Z8254: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_23,
    S => R1IN_ADD_2_1_AXB_24,
    LO => R1IN_ADD_2_1_CRY_24);
R1IN_ADD_2_1_S_23_Z8255: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_23,
    CI => R1IN_ADD_2_1_CRY_22,
    O => R1IN_ADD_2_1_S_23);
R1IN_ADD_2_1_CRY_23_Z8256: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_22,
    S => R1IN_ADD_2_1_AXB_23,
    LO => R1IN_ADD_2_1_CRY_23);
R1IN_ADD_2_1_S_22_Z8257: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_22,
    CI => R1IN_ADD_2_1_CRY_21,
    O => R1IN_ADD_2_1_S_22);
R1IN_ADD_2_1_CRY_22_Z8258: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_21,
    S => R1IN_ADD_2_1_AXB_22,
    LO => R1IN_ADD_2_1_CRY_22);
R1IN_ADD_2_1_S_21_Z8259: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_21,
    CI => R1IN_ADD_2_1_CRY_20,
    O => R1IN_ADD_2_1_S_21);
R1IN_ADD_2_1_CRY_21_Z8260: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_20,
    S => R1IN_ADD_2_1_AXB_21,
    LO => R1IN_ADD_2_1_CRY_21);
R1IN_ADD_2_1_S_20_Z8261: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_20,
    CI => R1IN_ADD_2_1_CRY_19,
    O => R1IN_ADD_2_1_S_20);
R1IN_ADD_2_1_CRY_20_Z8262: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_19,
    S => R1IN_ADD_2_1_AXB_20,
    LO => R1IN_ADD_2_1_CRY_20);
R1IN_ADD_2_1_S_19_Z8263: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_19,
    CI => R1IN_ADD_2_1_CRY_18,
    O => R1IN_ADD_2_1_S_19);
R1IN_ADD_2_1_CRY_19_Z8264: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_18,
    S => R1IN_ADD_2_1_AXB_19,
    LO => R1IN_ADD_2_1_CRY_19);
R1IN_ADD_2_1_S_18_Z8265: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_18,
    CI => R1IN_ADD_2_1_CRY_17,
    O => R1IN_ADD_2_1_S_18);
R1IN_ADD_2_1_CRY_18_Z8266: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_17,
    S => R1IN_ADD_2_1_AXB_18,
    LO => R1IN_ADD_2_1_CRY_18);
R1IN_ADD_2_1_S_17_Z8267: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_17,
    CI => R1IN_ADD_2_1_CRY_16,
    O => R1IN_ADD_2_1_S_17);
R1IN_ADD_2_1_CRY_17_Z8268: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_16,
    S => R1IN_ADD_2_1_AXB_17,
    LO => R1IN_ADD_2_1_CRY_17);
R1IN_ADD_2_1_S_16_Z8269: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_16,
    CI => R1IN_ADD_2_1_CRY_15,
    O => R1IN_ADD_2_1_S_16);
R1IN_ADD_2_1_CRY_16_Z8270: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_15,
    S => R1IN_ADD_2_1_AXB_16,
    LO => R1IN_ADD_2_1_CRY_16);
R1IN_ADD_2_1_S_15_Z8271: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_15,
    CI => R1IN_ADD_2_1_CRY_14,
    O => R1IN_ADD_2_1_S_15);
R1IN_ADD_2_1_CRY_15_Z8272: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_14,
    S => R1IN_ADD_2_1_AXB_15,
    LO => R1IN_ADD_2_1_CRY_15);
R1IN_ADD_2_1_S_14_Z8273: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_14,
    CI => R1IN_ADD_2_1_CRY_13,
    O => R1IN_ADD_2_1_S_14);
R1IN_ADD_2_1_CRY_14_Z8274: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_13,
    S => R1IN_ADD_2_1_AXB_14,
    LO => R1IN_ADD_2_1_CRY_14);
R1IN_ADD_2_1_S_13_Z8275: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_13,
    CI => R1IN_ADD_2_1_CRY_12,
    O => R1IN_ADD_2_1_S_13);
R1IN_ADD_2_1_CRY_13_Z8276: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_12,
    S => R1IN_ADD_2_1_AXB_13,
    LO => R1IN_ADD_2_1_CRY_13);
R1IN_ADD_2_1_S_12_Z8277: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_12,
    CI => R1IN_ADD_2_1_CRY_11,
    O => R1IN_ADD_2_1_S_12);
R1IN_ADD_2_1_CRY_12_Z8278: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_11,
    S => R1IN_ADD_2_1_AXB_12,
    LO => R1IN_ADD_2_1_CRY_12);
R1IN_ADD_2_1_S_11_Z8279: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_11,
    CI => R1IN_ADD_2_1_CRY_10,
    O => R1IN_ADD_2_1_S_11);
R1IN_ADD_2_1_CRY_11_Z8280: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_10,
    S => R1IN_ADD_2_1_AXB_11,
    LO => R1IN_ADD_2_1_CRY_11);
R1IN_ADD_2_1_S_10_Z8281: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_10,
    CI => R1IN_ADD_2_1_CRY_9,
    O => R1IN_ADD_2_1_S_10);
R1IN_ADD_2_1_CRY_10_Z8282: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_9,
    S => R1IN_ADD_2_1_AXB_10,
    LO => R1IN_ADD_2_1_CRY_10);
R1IN_ADD_2_1_S_9_Z8283: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_9,
    CI => R1IN_ADD_2_1_CRY_8,
    O => R1IN_ADD_2_1_S_9);
R1IN_ADD_2_1_CRY_9_Z8284: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_ADD_2_1_CRY_8,
    S => R1IN_ADD_2_1_AXB_9,
    LO => R1IN_ADD_2_1_CRY_9);
R1IN_ADD_2_1_S_8_Z8285: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_8,
    CI => R1IN_ADD_2_1_CRY_7,
    O => R1IN_ADD_2_1_S_8);
R1IN_ADD_2_1_CRY_8_Z8286: MUXCY_L port map (
    DI => R1IN_4F(44),
    CI => R1IN_ADD_2_1_CRY_7,
    S => R1IN_ADD_2_1_AXB_8,
    LO => R1IN_ADD_2_1_CRY_8);
R1IN_ADD_2_1_S_7_Z8287: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_7,
    CI => R1IN_ADD_2_1_CRY_6,
    O => R1IN_ADD_2_1_S_7);
R1IN_ADD_2_1_CRY_7_Z8288: MUXCY_L port map (
    DI => R1IN_4F(43),
    CI => R1IN_ADD_2_1_CRY_6,
    S => R1IN_ADD_2_1_AXB_7,
    LO => R1IN_ADD_2_1_CRY_7);
R1IN_ADD_2_1_S_6_Z8289: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_6,
    CI => R1IN_ADD_2_1_CRY_5,
    O => R1IN_ADD_2_1_S_6);
R1IN_ADD_2_1_CRY_6_Z8290: MUXCY_L port map (
    DI => R1IN_4F(42),
    CI => R1IN_ADD_2_1_CRY_5,
    S => R1IN_ADD_2_1_AXB_6,
    LO => R1IN_ADD_2_1_CRY_6);
R1IN_ADD_2_1_S_5_Z8291: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_5,
    CI => R1IN_ADD_2_1_CRY_4,
    O => R1IN_ADD_2_1_S_5);
R1IN_ADD_2_1_CRY_5_Z8292: MUXCY_L port map (
    DI => R1IN_4F(41),
    CI => R1IN_ADD_2_1_CRY_4,
    S => R1IN_ADD_2_1_AXB_5,
    LO => R1IN_ADD_2_1_CRY_5);
R1IN_ADD_2_1_S_4_Z8293: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_4,
    CI => R1IN_ADD_2_1_CRY_3,
    O => R1IN_ADD_2_1_S_4);
R1IN_ADD_2_1_CRY_4_Z8294: MUXCY_L port map (
    DI => R1IN_4F(40),
    CI => R1IN_ADD_2_1_CRY_3,
    S => R1IN_ADD_2_1_AXB_4,
    LO => R1IN_ADD_2_1_CRY_4);
R1IN_ADD_2_1_S_3_Z8295: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_3,
    CI => R1IN_ADD_2_1_CRY_2,
    O => R1IN_ADD_2_1_S_3);
R1IN_ADD_2_1_CRY_3_Z8296: MUXCY_L port map (
    DI => R1IN_4F(39),
    CI => R1IN_ADD_2_1_CRY_2,
    S => R1IN_ADD_2_1_AXB_3,
    LO => R1IN_ADD_2_1_CRY_3);
R1IN_ADD_2_1_S_2_Z8297: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_2,
    CI => R1IN_ADD_2_1_CRY_1,
    O => R1IN_ADD_2_1_S_2);
R1IN_ADD_2_1_CRY_2_Z8298: MUXCY_L port map (
    DI => R1IN_4F(38),
    CI => R1IN_ADD_2_1_CRY_1,
    S => R1IN_ADD_2_1_AXB_2,
    LO => R1IN_ADD_2_1_CRY_2);
R1IN_ADD_2_1_S_1_Z8299: XORCY port map (
    LI => R1IN_ADD_2_1_AXB_1,
    CI => R1IN_ADD_2_1_CRY_0,
    O => R1IN_ADD_2_1_S_1);
R1IN_ADD_2_1_CRY_1_Z8300: MUXCY_L port map (
    DI => R1IN_4F(37),
    CI => R1IN_ADD_2_1_CRY_0,
    S => R1IN_ADD_2_1_AXB_1,
    LO => R1IN_ADD_2_1_CRY_1);
R1IN_ADD_2_1_CRY_0_Z8301: MUXCY_L port map (
    DI => R1IN_4F(36),
    CI => NN_1,
    S => R1IN_ADD_2_1_AXB_0,
    LO => R1IN_ADD_2_1_CRY_0);
R1IN_ADD_2_0_S_52: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_52,
    CI => R1IN_ADD_2_0_CRY_51,
    O => PRODUCT(69));
R1IN_ADD_2_0_CRY_52_Z8303: MUXCY port map (
    DI => R1IN_4F(35),
    CI => R1IN_ADD_2_0_CRY_51,
    S => R1IN_ADD_2_0_AXB_52,
    O => R1IN_ADD_2_0_CRY_52);
R1IN_ADD_2_0_S_51: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_51,
    CI => R1IN_ADD_2_0_CRY_50,
    O => PRODUCT(68));
R1IN_ADD_2_0_CRY_51_Z8305: MUXCY_L port map (
    DI => R1IN_4F(34),
    CI => R1IN_ADD_2_0_CRY_50,
    S => R1IN_ADD_2_0_AXB_51,
    LO => R1IN_ADD_2_0_CRY_51);
R1IN_ADD_2_0_S_50: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_50,
    CI => R1IN_ADD_2_0_CRY_49,
    O => PRODUCT(67));
R1IN_ADD_2_0_CRY_50_Z8307: MUXCY_L port map (
    DI => R1IN_4F(33),
    CI => R1IN_ADD_2_0_CRY_49,
    S => R1IN_ADD_2_0_AXB_50,
    LO => R1IN_ADD_2_0_CRY_50);
R1IN_ADD_2_0_S_49: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_49,
    CI => R1IN_ADD_2_0_CRY_48,
    O => PRODUCT(66));
R1IN_ADD_2_0_CRY_49_Z8309: MUXCY_L port map (
    DI => R1IN_4F(32),
    CI => R1IN_ADD_2_0_CRY_48,
    S => R1IN_ADD_2_0_AXB_49,
    LO => R1IN_ADD_2_0_CRY_49);
R1IN_ADD_2_0_S_48: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_48,
    CI => R1IN_ADD_2_0_CRY_47,
    O => PRODUCT(65));
R1IN_ADD_2_0_CRY_48_Z8311: MUXCY_L port map (
    DI => R1IN_4F(31),
    CI => R1IN_ADD_2_0_CRY_47,
    S => R1IN_ADD_2_0_AXB_48,
    LO => R1IN_ADD_2_0_CRY_48);
R1IN_ADD_2_0_S_47: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_47,
    CI => R1IN_ADD_2_0_CRY_46,
    O => PRODUCT(64));
R1IN_ADD_2_0_CRY_47_Z8313: MUXCY_L port map (
    DI => R1IN_4F(30),
    CI => R1IN_ADD_2_0_CRY_46,
    S => R1IN_ADD_2_0_AXB_47,
    LO => R1IN_ADD_2_0_CRY_47);
R1IN_ADD_2_0_S_46: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_46,
    CI => R1IN_ADD_2_0_CRY_45,
    O => PRODUCT(63));
R1IN_ADD_2_0_CRY_46_Z8315: MUXCY_L port map (
    DI => R1IN_4F(29),
    CI => R1IN_ADD_2_0_CRY_45,
    S => R1IN_ADD_2_0_AXB_46,
    LO => R1IN_ADD_2_0_CRY_46);
R1IN_ADD_2_0_S_45: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_45,
    CI => R1IN_ADD_2_0_CRY_44,
    O => PRODUCT(62));
R1IN_ADD_2_0_CRY_45_Z8317: MUXCY_L port map (
    DI => R1IN_4F(28),
    CI => R1IN_ADD_2_0_CRY_44,
    S => R1IN_ADD_2_0_AXB_45,
    LO => R1IN_ADD_2_0_CRY_45);
R1IN_ADD_2_0_S_44: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_44,
    CI => R1IN_ADD_2_0_CRY_43,
    O => PRODUCT(61));
R1IN_ADD_2_0_CRY_44_Z8319: MUXCY_L port map (
    DI => R1IN_4F(27),
    CI => R1IN_ADD_2_0_CRY_43,
    S => R1IN_ADD_2_0_AXB_44,
    LO => R1IN_ADD_2_0_CRY_44);
R1IN_ADD_2_0_S_43: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_43,
    CI => R1IN_ADD_2_0_CRY_42,
    O => PRODUCT(60));
R1IN_ADD_2_0_CRY_43_Z8321: MUXCY_L port map (
    DI => R1IN_4F(26),
    CI => R1IN_ADD_2_0_CRY_42,
    S => R1IN_ADD_2_0_AXB_43,
    LO => R1IN_ADD_2_0_CRY_43);
R1IN_ADD_2_0_S_42: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_42,
    CI => R1IN_ADD_2_0_CRY_41,
    O => PRODUCT(59));
R1IN_ADD_2_0_CRY_42_Z8323: MUXCY_L port map (
    DI => R1IN_4F(25),
    CI => R1IN_ADD_2_0_CRY_41,
    S => R1IN_ADD_2_0_AXB_42,
    LO => R1IN_ADD_2_0_CRY_42);
R1IN_ADD_2_0_S_41: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_41,
    CI => R1IN_ADD_2_0_CRY_40,
    O => PRODUCT(58));
R1IN_ADD_2_0_CRY_41_Z8325: MUXCY_L port map (
    DI => R1IN_4F(24),
    CI => R1IN_ADD_2_0_CRY_40,
    S => R1IN_ADD_2_0_AXB_41,
    LO => R1IN_ADD_2_0_CRY_41);
R1IN_ADD_2_0_S_40: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_40,
    CI => R1IN_ADD_2_0_CRY_39,
    O => PRODUCT(57));
R1IN_ADD_2_0_CRY_40_Z8327: MUXCY_L port map (
    DI => R1IN_4F(23),
    CI => R1IN_ADD_2_0_CRY_39,
    S => R1IN_ADD_2_0_AXB_40,
    LO => R1IN_ADD_2_0_CRY_40);
R1IN_ADD_2_0_S_39: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_39,
    CI => R1IN_ADD_2_0_CRY_38,
    O => PRODUCT(56));
R1IN_ADD_2_0_CRY_39_Z8329: MUXCY_L port map (
    DI => R1IN_4F(22),
    CI => R1IN_ADD_2_0_CRY_38,
    S => R1IN_ADD_2_0_AXB_39,
    LO => R1IN_ADD_2_0_CRY_39);
R1IN_ADD_2_0_S_38: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_38,
    CI => R1IN_ADD_2_0_CRY_37,
    O => PRODUCT(55));
R1IN_ADD_2_0_CRY_38_Z8331: MUXCY_L port map (
    DI => R1IN_4F(21),
    CI => R1IN_ADD_2_0_CRY_37,
    S => R1IN_ADD_2_0_AXB_38,
    LO => R1IN_ADD_2_0_CRY_38);
R1IN_ADD_2_0_S_37: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_37,
    CI => R1IN_ADD_2_0_CRY_36,
    O => PRODUCT(54));
R1IN_ADD_2_0_CRY_37_Z8333: MUXCY_L port map (
    DI => R1IN_4F(20),
    CI => R1IN_ADD_2_0_CRY_36,
    S => R1IN_ADD_2_0_AXB_37,
    LO => R1IN_ADD_2_0_CRY_37);
R1IN_ADD_2_0_S_36: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_36,
    CI => R1IN_ADD_2_0_CRY_35,
    O => PRODUCT(53));
R1IN_ADD_2_0_CRY_36_Z8335: MUXCY_L port map (
    DI => R1IN_4F(19),
    CI => R1IN_ADD_2_0_CRY_35,
    S => R1IN_ADD_2_0_AXB_36,
    LO => R1IN_ADD_2_0_CRY_36);
R1IN_ADD_2_0_S_35: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_35,
    CI => R1IN_ADD_2_0_CRY_34,
    O => PRODUCT(52));
R1IN_ADD_2_0_CRY_35_Z8337: MUXCY_L port map (
    DI => R1IN_4F(18),
    CI => R1IN_ADD_2_0_CRY_34,
    S => R1IN_ADD_2_0_AXB_35,
    LO => R1IN_ADD_2_0_CRY_35);
R1IN_ADD_2_0_S_34: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_34,
    CI => R1IN_ADD_2_0_CRY_33,
    O => PRODUCT(51));
R1IN_ADD_2_0_CRY_34_Z8339: MUXCY_L port map (
    DI => R1IN_4F(17),
    CI => R1IN_ADD_2_0_CRY_33,
    S => R1IN_ADD_2_0_AXB_34,
    LO => R1IN_ADD_2_0_CRY_34);
R1IN_ADD_2_0_S_33: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_33,
    CI => R1IN_ADD_2_0_CRY_32,
    O => PRODUCT(50));
R1IN_ADD_2_0_CRY_33_Z8341: MUXCY_L port map (
    DI => R1IN_4FF(16),
    CI => R1IN_ADD_2_0_CRY_32,
    S => R1IN_ADD_2_0_AXB_33,
    LO => R1IN_ADD_2_0_CRY_33);
R1IN_ADD_2_0_S_32: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_32,
    CI => R1IN_ADD_2_0_CRY_31,
    O => PRODUCT(49));
R1IN_ADD_2_0_CRY_32_Z8343: MUXCY_L port map (
    DI => R1IN_4FF(15),
    CI => R1IN_ADD_2_0_CRY_31,
    S => R1IN_ADD_2_0_AXB_32,
    LO => R1IN_ADD_2_0_CRY_32);
R1IN_ADD_2_0_S_31: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_31,
    CI => R1IN_ADD_2_0_CRY_30,
    O => PRODUCT(48));
R1IN_ADD_2_0_CRY_31_Z8345: MUXCY_L port map (
    DI => R1IN_4FF(14),
    CI => R1IN_ADD_2_0_CRY_30,
    S => R1IN_ADD_2_0_AXB_31,
    LO => R1IN_ADD_2_0_CRY_31);
R1IN_ADD_2_0_S_30: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_30,
    CI => R1IN_ADD_2_0_CRY_29,
    O => PRODUCT(47));
R1IN_ADD_2_0_CRY_30_Z8347: MUXCY_L port map (
    DI => R1IN_4FF(13),
    CI => R1IN_ADD_2_0_CRY_29,
    S => R1IN_ADD_2_0_AXB_30,
    LO => R1IN_ADD_2_0_CRY_30);
R1IN_ADD_2_0_S_29: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_29,
    CI => R1IN_ADD_2_0_CRY_28,
    O => PRODUCT(46));
R1IN_ADD_2_0_CRY_29_Z8349: MUXCY_L port map (
    DI => R1IN_4FF(12),
    CI => R1IN_ADD_2_0_CRY_28,
    S => R1IN_ADD_2_0_AXB_29,
    LO => R1IN_ADD_2_0_CRY_29);
R1IN_ADD_2_0_S_28: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_28,
    CI => R1IN_ADD_2_0_CRY_27,
    O => PRODUCT(45));
R1IN_ADD_2_0_CRY_28_Z8351: MUXCY_L port map (
    DI => R1IN_4FF(11),
    CI => R1IN_ADD_2_0_CRY_27,
    S => R1IN_ADD_2_0_AXB_28,
    LO => R1IN_ADD_2_0_CRY_28);
R1IN_ADD_2_0_S_27: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_27,
    CI => R1IN_ADD_2_0_CRY_26,
    O => PRODUCT(44));
R1IN_ADD_2_0_CRY_27_Z8353: MUXCY_L port map (
    DI => R1IN_4FF(10),
    CI => R1IN_ADD_2_0_CRY_26,
    S => R1IN_ADD_2_0_AXB_27,
    LO => R1IN_ADD_2_0_CRY_27);
R1IN_ADD_2_0_S_26: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_26,
    CI => R1IN_ADD_2_0_CRY_25,
    O => PRODUCT(43));
R1IN_ADD_2_0_CRY_26_Z8355: MUXCY_L port map (
    DI => R1IN_4FF(9),
    CI => R1IN_ADD_2_0_CRY_25,
    S => R1IN_ADD_2_0_AXB_26,
    LO => R1IN_ADD_2_0_CRY_26);
R1IN_ADD_2_0_S_25: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_25,
    CI => R1IN_ADD_2_0_CRY_24,
    O => PRODUCT(42));
R1IN_ADD_2_0_CRY_25_Z8357: MUXCY_L port map (
    DI => R1IN_4FF(8),
    CI => R1IN_ADD_2_0_CRY_24,
    S => R1IN_ADD_2_0_AXB_25,
    LO => R1IN_ADD_2_0_CRY_25);
R1IN_ADD_2_0_S_24: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_24,
    CI => R1IN_ADD_2_0_CRY_23,
    O => PRODUCT(41));
R1IN_ADD_2_0_CRY_24_Z8359: MUXCY_L port map (
    DI => R1IN_4FF(7),
    CI => R1IN_ADD_2_0_CRY_23,
    S => R1IN_ADD_2_0_AXB_24,
    LO => R1IN_ADD_2_0_CRY_24);
R1IN_ADD_2_0_S_23: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_23,
    CI => R1IN_ADD_2_0_CRY_22,
    O => PRODUCT(40));
R1IN_ADD_2_0_CRY_23_Z8361: MUXCY_L port map (
    DI => R1IN_4FF(6),
    CI => R1IN_ADD_2_0_CRY_22,
    S => R1IN_ADD_2_0_AXB_23,
    LO => R1IN_ADD_2_0_CRY_23);
R1IN_ADD_2_0_S_22: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_22,
    CI => R1IN_ADD_2_0_CRY_21,
    O => PRODUCT(39));
R1IN_ADD_2_0_CRY_22_Z8363: MUXCY_L port map (
    DI => R1IN_4FF(5),
    CI => R1IN_ADD_2_0_CRY_21,
    S => R1IN_ADD_2_0_AXB_22,
    LO => R1IN_ADD_2_0_CRY_22);
R1IN_ADD_2_0_S_21: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_21,
    CI => R1IN_ADD_2_0_CRY_20,
    O => PRODUCT(38));
R1IN_ADD_2_0_CRY_21_Z8365: MUXCY_L port map (
    DI => R1IN_4FF(4),
    CI => R1IN_ADD_2_0_CRY_20,
    S => R1IN_ADD_2_0_AXB_21,
    LO => R1IN_ADD_2_0_CRY_21);
R1IN_ADD_2_0_S_20: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_20,
    CI => R1IN_ADD_2_0_CRY_19,
    O => PRODUCT(37));
R1IN_ADD_2_0_CRY_20_Z8367: MUXCY_L port map (
    DI => R1IN_4FF(3),
    CI => R1IN_ADD_2_0_CRY_19,
    S => R1IN_ADD_2_0_AXB_20,
    LO => R1IN_ADD_2_0_CRY_20);
R1IN_ADD_2_0_S_19: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_19,
    CI => R1IN_ADD_2_0_CRY_18,
    O => PRODUCT(36));
R1IN_ADD_2_0_CRY_19_Z8369: MUXCY_L port map (
    DI => R1IN_4FF(2),
    CI => R1IN_ADD_2_0_CRY_18,
    S => R1IN_ADD_2_0_AXB_19,
    LO => R1IN_ADD_2_0_CRY_19);
R1IN_ADD_2_0_S_18: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_18,
    CI => R1IN_ADD_2_0_CRY_17,
    O => PRODUCT(35));
R1IN_ADD_2_0_CRY_18_Z8371: MUXCY_L port map (
    DI => R1IN_4FF(1),
    CI => R1IN_ADD_2_0_CRY_17,
    S => R1IN_ADD_2_0_AXB_18,
    LO => R1IN_ADD_2_0_CRY_18);
R1IN_ADD_2_0_S_17: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_17,
    CI => R1IN_ADD_2_0_CRY_16,
    O => PRODUCT(34));
R1IN_ADD_2_0_CRY_17_Z8373: MUXCY_L port map (
    DI => R1IN_4FF(0),
    CI => R1IN_ADD_2_0_CRY_16,
    S => R1IN_ADD_2_0_AXB_17,
    LO => R1IN_ADD_2_0_CRY_17);
R1IN_ADD_2_0_S_16: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_16,
    CI => R1IN_ADD_2_0_CRY_15,
    O => PRODUCT(33));
R1IN_ADD_2_0_CRY_16_Z8375: MUXCY_L port map (
    DI => R1IN_1FF(33),
    CI => R1IN_ADD_2_0_CRY_15,
    S => R1IN_ADD_2_0_AXB_16,
    LO => R1IN_ADD_2_0_CRY_16);
R1IN_ADD_2_0_S_15: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_15,
    CI => R1IN_ADD_2_0_CRY_14,
    O => PRODUCT(32));
R1IN_ADD_2_0_CRY_15_Z8377: MUXCY_L port map (
    DI => R1IN_1FF(32),
    CI => R1IN_ADD_2_0_CRY_14,
    S => R1IN_ADD_2_0_AXB_15,
    LO => R1IN_ADD_2_0_CRY_15);
R1IN_ADD_2_0_S_14: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_14,
    CI => R1IN_ADD_2_0_CRY_13,
    O => PRODUCT(31));
R1IN_ADD_2_0_CRY_14_Z8379: MUXCY_L port map (
    DI => R1IN_1FF(31),
    CI => R1IN_ADD_2_0_CRY_13,
    S => R1IN_ADD_2_0_AXB_14,
    LO => R1IN_ADD_2_0_CRY_14);
R1IN_ADD_2_0_S_13: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_13,
    CI => R1IN_ADD_2_0_CRY_12,
    O => PRODUCT(30));
R1IN_ADD_2_0_CRY_13_Z8381: MUXCY_L port map (
    DI => R1IN_1FF(30),
    CI => R1IN_ADD_2_0_CRY_12,
    S => R1IN_ADD_2_0_AXB_13,
    LO => R1IN_ADD_2_0_CRY_13);
R1IN_ADD_2_0_S_12: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_12,
    CI => R1IN_ADD_2_0_CRY_11,
    O => PRODUCT(29));
R1IN_ADD_2_0_CRY_12_Z8383: MUXCY_L port map (
    DI => R1IN_1FF(29),
    CI => R1IN_ADD_2_0_CRY_11,
    S => R1IN_ADD_2_0_AXB_12,
    LO => R1IN_ADD_2_0_CRY_12);
R1IN_ADD_2_0_S_11: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_11,
    CI => R1IN_ADD_2_0_CRY_10,
    O => PRODUCT(28));
R1IN_ADD_2_0_CRY_11_Z8385: MUXCY_L port map (
    DI => R1IN_1FF(28),
    CI => R1IN_ADD_2_0_CRY_10,
    S => R1IN_ADD_2_0_AXB_11,
    LO => R1IN_ADD_2_0_CRY_11);
R1IN_ADD_2_0_S_10: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_10,
    CI => R1IN_ADD_2_0_CRY_9,
    O => PRODUCT(27));
R1IN_ADD_2_0_CRY_10_Z8387: MUXCY_L port map (
    DI => R1IN_1FF(27),
    CI => R1IN_ADD_2_0_CRY_9,
    S => R1IN_ADD_2_0_AXB_10,
    LO => R1IN_ADD_2_0_CRY_10);
R1IN_ADD_2_0_S_9: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_9,
    CI => R1IN_ADD_2_0_CRY_8,
    O => PRODUCT(26));
R1IN_ADD_2_0_CRY_9_Z8389: MUXCY_L port map (
    DI => R1IN_1FF(26),
    CI => R1IN_ADD_2_0_CRY_8,
    S => R1IN_ADD_2_0_AXB_9,
    LO => R1IN_ADD_2_0_CRY_9);
R1IN_ADD_2_0_S_8: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_8,
    CI => R1IN_ADD_2_0_CRY_7,
    O => PRODUCT(25));
R1IN_ADD_2_0_CRY_8_Z8391: MUXCY_L port map (
    DI => R1IN_1FF(25),
    CI => R1IN_ADD_2_0_CRY_7,
    S => R1IN_ADD_2_0_AXB_8,
    LO => R1IN_ADD_2_0_CRY_8);
R1IN_ADD_2_0_S_7: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_7,
    CI => R1IN_ADD_2_0_CRY_6,
    O => PRODUCT(24));
R1IN_ADD_2_0_CRY_7_Z8393: MUXCY_L port map (
    DI => R1IN_1FF(24),
    CI => R1IN_ADD_2_0_CRY_6,
    S => R1IN_ADD_2_0_AXB_7,
    LO => R1IN_ADD_2_0_CRY_7);
R1IN_ADD_2_0_S_6: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_6,
    CI => R1IN_ADD_2_0_CRY_5,
    O => PRODUCT(23));
R1IN_ADD_2_0_CRY_6_Z8395: MUXCY_L port map (
    DI => R1IN_1FF(23),
    CI => R1IN_ADD_2_0_CRY_5,
    S => R1IN_ADD_2_0_AXB_6,
    LO => R1IN_ADD_2_0_CRY_6);
R1IN_ADD_2_0_S_5: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_5,
    CI => R1IN_ADD_2_0_CRY_4,
    O => PRODUCT(22));
R1IN_ADD_2_0_CRY_5_Z8397: MUXCY_L port map (
    DI => R1IN_1FF(22),
    CI => R1IN_ADD_2_0_CRY_4,
    S => R1IN_ADD_2_0_AXB_5,
    LO => R1IN_ADD_2_0_CRY_5);
R1IN_ADD_2_0_S_4: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_4,
    CI => R1IN_ADD_2_0_CRY_3,
    O => PRODUCT(21));
R1IN_ADD_2_0_CRY_4_Z8399: MUXCY_L port map (
    DI => R1IN_1FF(21),
    CI => R1IN_ADD_2_0_CRY_3,
    S => R1IN_ADD_2_0_AXB_4,
    LO => R1IN_ADD_2_0_CRY_4);
R1IN_ADD_2_0_S_3: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_3,
    CI => R1IN_ADD_2_0_CRY_2,
    O => PRODUCT(20));
R1IN_ADD_2_0_CRY_3_Z8401: MUXCY_L port map (
    DI => R1IN_1FF(20),
    CI => R1IN_ADD_2_0_CRY_2,
    S => R1IN_ADD_2_0_AXB_3,
    LO => R1IN_ADD_2_0_CRY_3);
R1IN_ADD_2_0_S_2: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_2,
    CI => R1IN_ADD_2_0_CRY_1,
    O => PRODUCT(19));
R1IN_ADD_2_0_CRY_2_Z8403: MUXCY_L port map (
    DI => R1IN_1FF(19),
    CI => R1IN_ADD_2_0_CRY_1,
    S => R1IN_ADD_2_0_AXB_2,
    LO => R1IN_ADD_2_0_CRY_2);
R1IN_ADD_2_0_S_1: XORCY port map (
    LI => R1IN_ADD_2_0_AXB_1,
    CI => R1IN_ADD_2_0_CRY_0,
    O => PRODUCT(18));
R1IN_ADD_2_0_CRY_1_Z8405: MUXCY_L port map (
    DI => R1IN_1FF(18),
    CI => R1IN_ADD_2_0_CRY_0,
    S => R1IN_ADD_2_0_AXB_1,
    LO => R1IN_ADD_2_0_CRY_1);
R1IN_ADD_2_0_CRY_0_Z8406: MUXCY_L port map (
    DI => R1IN_ADD_2_0,
    CI => NN_1,
    S => NN_11,
    LO => R1IN_ADD_2_0_CRY_0);
R1IN_4_ADD_2_1_S_34: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_34,
    CI => R1IN_4_ADD_2_1_CRY_33,
    O => N_1781_RETI);
R1IN_4_ADD_2_1_S_33: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_33,
    CI => R1IN_4_ADD_2_1_CRY_32,
    O => N_1779_RETI);
R1IN_4_ADD_2_1_CRY_33_Z8409: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_32,
    S => R1IN_4_ADD_2_1_AXB_33,
    LO => R1IN_4_ADD_2_1_CRY_33);
R1IN_4_ADD_2_1_S_32: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_32,
    CI => R1IN_4_ADD_2_1_CRY_31,
    O => N_1777_RETI);
R1IN_4_ADD_2_1_CRY_32_Z8411: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_31,
    S => R1IN_4_ADD_2_1_AXB_32,
    LO => R1IN_4_ADD_2_1_CRY_32);
R1IN_4_ADD_2_1_S_31: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_31,
    CI => R1IN_4_ADD_2_1_CRY_30,
    O => N_1775_RETI);
R1IN_4_ADD_2_1_CRY_31_Z8413: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_30,
    S => R1IN_4_ADD_2_1_AXB_31,
    LO => R1IN_4_ADD_2_1_CRY_31);
R1IN_4_ADD_2_1_S_30: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_30,
    CI => R1IN_4_ADD_2_1_CRY_29,
    O => N_1773_RETI);
R1IN_4_ADD_2_1_CRY_30_Z8415: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_29,
    S => R1IN_4_ADD_2_1_AXB_30,
    LO => R1IN_4_ADD_2_1_CRY_30);
R1IN_4_ADD_2_1_S_29: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_29,
    CI => R1IN_4_ADD_2_1_CRY_28,
    O => N_1771_RETI);
R1IN_4_ADD_2_1_CRY_29_Z8417: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_28,
    S => R1IN_4_ADD_2_1_AXB_29,
    LO => R1IN_4_ADD_2_1_CRY_29);
R1IN_4_ADD_2_1_S_28: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_28,
    CI => R1IN_4_ADD_2_1_CRY_27,
    O => N_1769_RETI);
R1IN_4_ADD_2_1_CRY_28_Z8419: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_27,
    S => R1IN_4_ADD_2_1_AXB_28,
    LO => R1IN_4_ADD_2_1_CRY_28);
R1IN_4_ADD_2_1_S_27: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_27,
    CI => R1IN_4_ADD_2_1_CRY_26,
    O => N_1767_RETI);
R1IN_4_ADD_2_1_CRY_27_Z8421: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_26,
    S => R1IN_4_ADD_2_1_AXB_27,
    LO => R1IN_4_ADD_2_1_CRY_27);
R1IN_4_ADD_2_1_S_26: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_26,
    CI => R1IN_4_ADD_2_1_CRY_25,
    O => N_1765_RETI);
R1IN_4_ADD_2_1_CRY_26_Z8423: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_25,
    S => R1IN_4_ADD_2_1_AXB_26,
    LO => R1IN_4_ADD_2_1_CRY_26);
R1IN_4_ADD_2_1_S_25: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_25,
    CI => R1IN_4_ADD_2_1_CRY_24,
    O => N_1763_RETI);
R1IN_4_ADD_2_1_CRY_25_Z8425: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_24,
    S => R1IN_4_ADD_2_1_AXB_25,
    LO => R1IN_4_ADD_2_1_CRY_25);
R1IN_4_ADD_2_1_S_24: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_24,
    CI => R1IN_4_ADD_2_1_CRY_23,
    O => N_1761_RETI);
R1IN_4_ADD_2_1_CRY_24_Z8427: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_23,
    S => R1IN_4_ADD_2_1_AXB_24,
    LO => R1IN_4_ADD_2_1_CRY_24);
R1IN_4_ADD_2_1_S_23: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_23,
    CI => R1IN_4_ADD_2_1_CRY_22,
    O => N_1759_RETI);
R1IN_4_ADD_2_1_CRY_23_Z8429: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_22,
    S => R1IN_4_ADD_2_1_AXB_23,
    LO => R1IN_4_ADD_2_1_CRY_23);
R1IN_4_ADD_2_1_S_22: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_22,
    CI => R1IN_4_ADD_2_1_CRY_21,
    O => N_1757_RETI);
R1IN_4_ADD_2_1_CRY_22_Z8431: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_21,
    S => R1IN_4_ADD_2_1_AXB_22,
    LO => R1IN_4_ADD_2_1_CRY_22);
R1IN_4_ADD_2_1_S_21: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_21,
    CI => R1IN_4_ADD_2_1_CRY_20,
    O => N_1755_RETI);
R1IN_4_ADD_2_1_CRY_21_Z8433: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_20,
    S => R1IN_4_ADD_2_1_AXB_21,
    LO => R1IN_4_ADD_2_1_CRY_21);
R1IN_4_ADD_2_1_S_20: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_20,
    CI => R1IN_4_ADD_2_1_CRY_19,
    O => N_1753_RETI);
R1IN_4_ADD_2_1_CRY_20_Z8435: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_19,
    S => R1IN_4_ADD_2_1_AXB_20,
    LO => R1IN_4_ADD_2_1_CRY_20);
R1IN_4_ADD_2_1_S_19: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_19,
    CI => R1IN_4_ADD_2_1_CRY_18,
    O => N_1751_RETI);
R1IN_4_ADD_2_1_CRY_19_Z8437: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_18,
    S => R1IN_4_ADD_2_1_AXB_19,
    LO => R1IN_4_ADD_2_1_CRY_19);
R1IN_4_ADD_2_1_S_18: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_18,
    CI => R1IN_4_ADD_2_1_CRY_17,
    O => N_1749_RETI);
R1IN_4_ADD_2_1_CRY_18_Z8439: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_17,
    S => R1IN_4_ADD_2_1_AXB_18,
    LO => R1IN_4_ADD_2_1_CRY_18);
R1IN_4_ADD_2_1_S_17: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_17,
    CI => R1IN_4_ADD_2_1_CRY_16,
    O => N_1747_RETI);
R1IN_4_ADD_2_1_CRY_17_Z8441: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_16,
    S => R1IN_4_ADD_2_1_AXB_17,
    LO => R1IN_4_ADD_2_1_CRY_17);
R1IN_4_ADD_2_1_S_16: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_16,
    CI => R1IN_4_ADD_2_1_CRY_15,
    O => N_1745_RETI);
R1IN_4_ADD_2_1_CRY_16_Z8443: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_15,
    S => R1IN_4_ADD_2_1_AXB_16,
    LO => R1IN_4_ADD_2_1_CRY_16);
R1IN_4_ADD_2_1_S_15: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_15,
    CI => R1IN_4_ADD_2_1_CRY_14,
    O => N_1743_RETI);
R1IN_4_ADD_2_1_CRY_15_Z8445: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_14,
    S => R1IN_4_ADD_2_1_AXB_15,
    LO => R1IN_4_ADD_2_1_CRY_15);
R1IN_4_ADD_2_1_S_14: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_14,
    CI => R1IN_4_ADD_2_1_CRY_13,
    O => N_1741_RETI);
R1IN_4_ADD_2_1_CRY_14_Z8447: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_13,
    S => R1IN_4_ADD_2_1_AXB_14,
    LO => R1IN_4_ADD_2_1_CRY_14);
R1IN_4_ADD_2_1_S_13: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_13,
    CI => R1IN_4_ADD_2_1_CRY_12,
    O => N_1739_RETI);
R1IN_4_ADD_2_1_CRY_13_Z8449: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_12,
    S => R1IN_4_ADD_2_1_AXB_13,
    LO => R1IN_4_ADD_2_1_CRY_13);
R1IN_4_ADD_2_1_S_12: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_12,
    CI => R1IN_4_ADD_2_1_CRY_11,
    O => N_1737_RETI);
R1IN_4_ADD_2_1_CRY_12_Z8451: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_11,
    S => R1IN_4_ADD_2_1_AXB_12,
    LO => R1IN_4_ADD_2_1_CRY_12);
R1IN_4_ADD_2_1_S_11: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_11,
    CI => R1IN_4_ADD_2_1_CRY_10,
    O => N_1735_RETI);
R1IN_4_ADD_2_1_CRY_11_Z8453: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_10,
    S => R1IN_4_ADD_2_1_AXB_11,
    LO => R1IN_4_ADD_2_1_CRY_11);
R1IN_4_ADD_2_1_S_10: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_10,
    CI => R1IN_4_ADD_2_1_CRY_9,
    O => N_1733_RETI);
R1IN_4_ADD_2_1_CRY_10_Z8455: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_9,
    S => R1IN_4_ADD_2_1_AXB_10,
    LO => R1IN_4_ADD_2_1_CRY_10);
R1IN_4_ADD_2_1_S_9: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_9,
    CI => R1IN_4_ADD_2_1_CRY_8,
    O => N_1731_RETI);
R1IN_4_ADD_2_1_CRY_9_Z8457: MUXCY_L port map (
    DI => NN_1,
    CI => R1IN_4_ADD_2_1_CRY_8,
    S => R1IN_4_ADD_2_1_AXB_9,
    LO => R1IN_4_ADD_2_1_CRY_9);
R1IN_4_ADD_2_1_S_8: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_8,
    CI => R1IN_4_ADD_2_1_CRY_7,
    O => N_1729_RETI);
R1IN_4_ADD_2_1_CRY_8_Z8459: MUXCY_L port map (
    DI => NN_10,
    CI => R1IN_4_ADD_2_1_CRY_7,
    S => R1IN_4_ADD_2_1_AXB_8,
    LO => R1IN_4_ADD_2_1_CRY_8);
R1IN_4_ADD_2_1_S_7: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_7,
    CI => R1IN_4_ADD_2_1_CRY_6,
    O => N_1727_RETI);
R1IN_4_ADD_2_1_CRY_7_Z8461: MUXCY_L port map (
    DI => NN_9,
    CI => R1IN_4_ADD_2_1_CRY_6,
    S => R1IN_4_ADD_2_1_AXB_7,
    LO => R1IN_4_ADD_2_1_CRY_7);
R1IN_4_ADD_2_1_S_6: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_6,
    CI => R1IN_4_ADD_2_1_CRY_5,
    O => N_1725_RETI);
R1IN_4_ADD_2_1_CRY_6_Z8463: MUXCY_L port map (
    DI => NN_8,
    CI => R1IN_4_ADD_2_1_CRY_5,
    S => R1IN_4_ADD_2_1_AXB_6,
    LO => R1IN_4_ADD_2_1_CRY_6);
R1IN_4_ADD_2_1_S_5: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_5,
    CI => R1IN_4_ADD_2_1_CRY_4,
    O => N_1723_RETI);
R1IN_4_ADD_2_1_CRY_5_Z8465: MUXCY_L port map (
    DI => NN_7,
    CI => R1IN_4_ADD_2_1_CRY_4,
    S => R1IN_4_ADD_2_1_AXB_5,
    LO => R1IN_4_ADD_2_1_CRY_5);
R1IN_4_ADD_2_1_S_4: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_4,
    CI => R1IN_4_ADD_2_1_CRY_3,
    O => N_1721_RETI);
R1IN_4_ADD_2_1_CRY_4_Z8467: MUXCY_L port map (
    DI => NN_6,
    CI => R1IN_4_ADD_2_1_CRY_3,
    S => R1IN_4_ADD_2_1_AXB_4,
    LO => R1IN_4_ADD_2_1_CRY_4);
R1IN_4_ADD_2_1_S_3: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_3,
    CI => R1IN_4_ADD_2_1_CRY_2,
    O => N_1719_RETI);
R1IN_4_ADD_2_1_CRY_3_Z8469: MUXCY_L port map (
    DI => NN_5,
    CI => R1IN_4_ADD_2_1_CRY_2,
    S => R1IN_4_ADD_2_1_AXB_3,
    LO => R1IN_4_ADD_2_1_CRY_3);
R1IN_4_ADD_2_1_S_2: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_2,
    CI => R1IN_4_ADD_2_1_CRY_1,
    O => N_1717_RETI);
R1IN_4_ADD_2_1_CRY_2_Z8471: MUXCY_L port map (
    DI => NN_4,
    CI => R1IN_4_ADD_2_1_CRY_1,
    S => R1IN_4_ADD_2_1_AXB_2,
    LO => R1IN_4_ADD_2_1_CRY_2);
R1IN_4_ADD_2_1_S_1: XORCY port map (
    LI => R1IN_4_ADD_2_1_AXB_1,
    CI => R1IN_4_ADD_2_1_CRY_0,
    O => N_1715_RETI);
R1IN_4_ADD_2_1_CRY_1_Z8473: MUXCY_L port map (
    DI => NN_3,
    CI => R1IN_4_ADD_2_1_CRY_0,
    S => R1IN_4_ADD_2_1_AXB_1,
    LO => R1IN_4_ADD_2_1_CRY_1);
R1IN_4_ADD_2_1_CRY_0_Z8474: MUXCY_L port map (
    DI => R1IN_4_ADD_2_1,
    CI => NN_1,
    S => R1IN_4_ADD_2_1_AXB_0_RETI,
    LO => R1IN_4_ADD_2_1_CRY_0);
R1IN_4_ADD_2_0_S_35: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_35,
    CI => R1IN_4_ADD_2_0_CRY_34,
    O => R1IN_4(52));
R1IN_4_ADD_2_0_CRY_35_Z8476: MUXCY port map (
    DI => R1IN_4_ADD_1(35),
    CI => R1IN_4_ADD_2_0_CRY_34,
    S => R1IN_4_ADD_2_0_AXB_35,
    O => R1IN_4_ADD_2_0_CRY_35);
R1IN_4_ADD_2_0_S_34: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_34,
    CI => R1IN_4_ADD_2_0_CRY_33,
    O => R1IN_4(51));
R1IN_4_ADD_2_0_CRY_34_Z8478: MUXCY_L port map (
    DI => R1IN_4_ADD_1(34),
    CI => R1IN_4_ADD_2_0_CRY_33,
    S => R1IN_4_ADD_2_0_AXB_34,
    LO => R1IN_4_ADD_2_0_CRY_34);
R1IN_4_ADD_2_0_S_33: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_33,
    CI => R1IN_4_ADD_2_0_CRY_32,
    O => R1IN_4(50));
R1IN_4_ADD_2_0_CRY_33_Z8480: MUXCY_L port map (
    DI => R1IN_4_ADD_1(33),
    CI => R1IN_4_ADD_2_0_CRY_32,
    S => R1IN_4_ADD_2_0_AXB_33,
    LO => R1IN_4_ADD_2_0_CRY_33);
R1IN_4_ADD_2_0_S_32: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_32,
    CI => R1IN_4_ADD_2_0_CRY_31,
    O => R1IN_4(49));
R1IN_4_ADD_2_0_CRY_32_Z8482: MUXCY_L port map (
    DI => R1IN_4_ADD_1(32),
    CI => R1IN_4_ADD_2_0_CRY_31,
    S => R1IN_4_ADD_2_0_AXB_32,
    LO => R1IN_4_ADD_2_0_CRY_32);
R1IN_4_ADD_2_0_S_31: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_31,
    CI => R1IN_4_ADD_2_0_CRY_30,
    O => R1IN_4(48));
R1IN_4_ADD_2_0_CRY_31_Z8484: MUXCY_L port map (
    DI => R1IN_4_ADD_1(31),
    CI => R1IN_4_ADD_2_0_CRY_30,
    S => R1IN_4_ADD_2_0_AXB_31,
    LO => R1IN_4_ADD_2_0_CRY_31);
R1IN_4_ADD_2_0_S_30: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_30,
    CI => R1IN_4_ADD_2_0_CRY_29,
    O => R1IN_4(47));
R1IN_4_ADD_2_0_CRY_30_Z8486: MUXCY_L port map (
    DI => R1IN_4_ADD_1(30),
    CI => R1IN_4_ADD_2_0_CRY_29,
    S => R1IN_4_ADD_2_0_AXB_30,
    LO => R1IN_4_ADD_2_0_CRY_30);
R1IN_4_ADD_2_0_S_29: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_29,
    CI => R1IN_4_ADD_2_0_CRY_28,
    O => R1IN_4(46));
R1IN_4_ADD_2_0_CRY_29_Z8488: MUXCY_L port map (
    DI => R1IN_4_ADD_1(29),
    CI => R1IN_4_ADD_2_0_CRY_28,
    S => R1IN_4_ADD_2_0_AXB_29,
    LO => R1IN_4_ADD_2_0_CRY_29);
R1IN_4_ADD_2_0_S_28: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_28,
    CI => R1IN_4_ADD_2_0_CRY_27,
    O => R1IN_4(45));
R1IN_4_ADD_2_0_CRY_28_Z8490: MUXCY_L port map (
    DI => R1IN_4_ADD_1(28),
    CI => R1IN_4_ADD_2_0_CRY_27,
    S => R1IN_4_ADD_2_0_AXB_28,
    LO => R1IN_4_ADD_2_0_CRY_28);
R1IN_4_ADD_2_0_S_27: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_27,
    CI => R1IN_4_ADD_2_0_CRY_26,
    O => R1IN_4(44));
R1IN_4_ADD_2_0_CRY_27_Z8492: MUXCY_L port map (
    DI => R1IN_4_ADD_1(27),
    CI => R1IN_4_ADD_2_0_CRY_26,
    S => R1IN_4_ADD_2_0_AXB_27,
    LO => R1IN_4_ADD_2_0_CRY_27);
R1IN_4_ADD_2_0_S_26: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_26,
    CI => R1IN_4_ADD_2_0_CRY_25,
    O => R1IN_4(43));
R1IN_4_ADD_2_0_CRY_26_Z8494: MUXCY_L port map (
    DI => R1IN_4_ADD_1(26),
    CI => R1IN_4_ADD_2_0_CRY_25,
    S => R1IN_4_ADD_2_0_AXB_26,
    LO => R1IN_4_ADD_2_0_CRY_26);
R1IN_4_ADD_2_0_S_25: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_25,
    CI => R1IN_4_ADD_2_0_CRY_24,
    O => R1IN_4(42));
R1IN_4_ADD_2_0_CRY_25_Z8496: MUXCY_L port map (
    DI => R1IN_4_ADD_1(25),
    CI => R1IN_4_ADD_2_0_CRY_24,
    S => R1IN_4_ADD_2_0_AXB_25,
    LO => R1IN_4_ADD_2_0_CRY_25);
R1IN_4_ADD_2_0_S_24: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_24,
    CI => R1IN_4_ADD_2_0_CRY_23,
    O => R1IN_4(41));
R1IN_4_ADD_2_0_CRY_24_Z8498: MUXCY_L port map (
    DI => R1IN_4_ADD_1(24),
    CI => R1IN_4_ADD_2_0_CRY_23,
    S => R1IN_4_ADD_2_0_AXB_24,
    LO => R1IN_4_ADD_2_0_CRY_24);
R1IN_4_ADD_2_0_S_23: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_23,
    CI => R1IN_4_ADD_2_0_CRY_22,
    O => R1IN_4(40));
R1IN_4_ADD_2_0_CRY_23_Z8500: MUXCY_L port map (
    DI => R1IN_4_ADD_1(23),
    CI => R1IN_4_ADD_2_0_CRY_22,
    S => R1IN_4_ADD_2_0_AXB_23,
    LO => R1IN_4_ADD_2_0_CRY_23);
R1IN_4_ADD_2_0_S_22: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_22,
    CI => R1IN_4_ADD_2_0_CRY_21,
    O => R1IN_4(39));
R1IN_4_ADD_2_0_CRY_22_Z8502: MUXCY_L port map (
    DI => R1IN_4_ADD_1(22),
    CI => R1IN_4_ADD_2_0_CRY_21,
    S => R1IN_4_ADD_2_0_AXB_22,
    LO => R1IN_4_ADD_2_0_CRY_22);
R1IN_4_ADD_2_0_S_21: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_21,
    CI => R1IN_4_ADD_2_0_CRY_20,
    O => R1IN_4(38));
R1IN_4_ADD_2_0_CRY_21_Z8504: MUXCY_L port map (
    DI => R1IN_4_ADD_1(21),
    CI => R1IN_4_ADD_2_0_CRY_20,
    S => R1IN_4_ADD_2_0_AXB_21,
    LO => R1IN_4_ADD_2_0_CRY_21);
R1IN_4_ADD_2_0_S_20: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_20,
    CI => R1IN_4_ADD_2_0_CRY_19,
    O => R1IN_4(37));
R1IN_4_ADD_2_0_CRY_20_Z8506: MUXCY_L port map (
    DI => R1IN_4_ADD_1(20),
    CI => R1IN_4_ADD_2_0_CRY_19,
    S => R1IN_4_ADD_2_0_AXB_20,
    LO => R1IN_4_ADD_2_0_CRY_20);
R1IN_4_ADD_2_0_S_19: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_19,
    CI => R1IN_4_ADD_2_0_CRY_18,
    O => R1IN_4(36));
R1IN_4_ADD_2_0_CRY_19_Z8508: MUXCY_L port map (
    DI => R1IN_4_ADD_1(19),
    CI => R1IN_4_ADD_2_0_CRY_18,
    S => R1IN_4_ADD_2_0_AXB_19,
    LO => R1IN_4_ADD_2_0_CRY_19);
R1IN_4_ADD_2_0_S_18: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_18,
    CI => R1IN_4_ADD_2_0_CRY_17,
    O => R1IN_4(35));
R1IN_4_ADD_2_0_CRY_18_Z8510: MUXCY_L port map (
    DI => R1IN_4_ADD_1(18),
    CI => R1IN_4_ADD_2_0_CRY_17,
    S => R1IN_4_ADD_2_0_AXB_18,
    LO => R1IN_4_ADD_2_0_CRY_18);
R1IN_4_ADD_2_0_S_17: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_17,
    CI => R1IN_4_ADD_2_0_CRY_16,
    O => R1IN_4(34));
R1IN_4_ADD_2_0_CRY_17_Z8512: MUXCY_L port map (
    DI => R1IN_4_ADD_1(17),
    CI => R1IN_4_ADD_2_0_CRY_16,
    S => R1IN_4_ADD_2_0_AXB_17,
    LO => R1IN_4_ADD_2_0_CRY_17);
R1IN_4_ADD_2_0_S_16: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_16,
    CI => R1IN_4_ADD_2_0_CRY_15,
    O => R1IN_4(33));
R1IN_4_ADD_2_0_CRY_16_Z8514: MUXCY_L port map (
    DI => R1IN_4_ADD_1(16),
    CI => R1IN_4_ADD_2_0_CRY_15,
    S => R1IN_4_ADD_2_0_AXB_16,
    LO => R1IN_4_ADD_2_0_CRY_16);
R1IN_4_ADD_2_0_S_15: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_15,
    CI => R1IN_4_ADD_2_0_CRY_14,
    O => R1IN_4(32));
R1IN_4_ADD_2_0_CRY_15_Z8516: MUXCY_L port map (
    DI => R1IN_4_ADD_1(15),
    CI => R1IN_4_ADD_2_0_CRY_14,
    S => R1IN_4_ADD_2_0_AXB_15,
    LO => R1IN_4_ADD_2_0_CRY_15);
R1IN_4_ADD_2_0_S_14: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_14,
    CI => R1IN_4_ADD_2_0_CRY_13,
    O => R1IN_4(31));
R1IN_4_ADD_2_0_CRY_14_Z8518: MUXCY_L port map (
    DI => R1IN_4_ADD_1(14),
    CI => R1IN_4_ADD_2_0_CRY_13,
    S => R1IN_4_ADD_2_0_AXB_14,
    LO => R1IN_4_ADD_2_0_CRY_14);
R1IN_4_ADD_2_0_S_13: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_13,
    CI => R1IN_4_ADD_2_0_CRY_12,
    O => R1IN_4(30));
R1IN_4_ADD_2_0_CRY_13_Z8520: MUXCY_L port map (
    DI => R1IN_4_ADD_1(13),
    CI => R1IN_4_ADD_2_0_CRY_12,
    S => R1IN_4_ADD_2_0_AXB_13,
    LO => R1IN_4_ADD_2_0_CRY_13);
R1IN_4_ADD_2_0_S_12: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_12,
    CI => R1IN_4_ADD_2_0_CRY_11,
    O => R1IN_4(29));
R1IN_4_ADD_2_0_CRY_12_Z8522: MUXCY_L port map (
    DI => R1IN_4_ADD_1(12),
    CI => R1IN_4_ADD_2_0_CRY_11,
    S => R1IN_4_ADD_2_0_AXB_12,
    LO => R1IN_4_ADD_2_0_CRY_12);
R1IN_4_ADD_2_0_S_11: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_11,
    CI => R1IN_4_ADD_2_0_CRY_10,
    O => R1IN_4(28));
R1IN_4_ADD_2_0_CRY_11_Z8524: MUXCY_L port map (
    DI => R1IN_4_ADD_1(11),
    CI => R1IN_4_ADD_2_0_CRY_10,
    S => R1IN_4_ADD_2_0_AXB_11,
    LO => R1IN_4_ADD_2_0_CRY_11);
R1IN_4_ADD_2_0_S_10: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_10,
    CI => R1IN_4_ADD_2_0_CRY_9,
    O => R1IN_4(27));
R1IN_4_ADD_2_0_CRY_10_Z8526: MUXCY_L port map (
    DI => R1IN_4_ADD_1(10),
    CI => R1IN_4_ADD_2_0_CRY_9,
    S => R1IN_4_ADD_2_0_AXB_10,
    LO => R1IN_4_ADD_2_0_CRY_10);
R1IN_4_ADD_2_0_S_9: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_9,
    CI => R1IN_4_ADD_2_0_CRY_8,
    O => R1IN_4(26));
R1IN_4_ADD_2_0_CRY_9_Z8528: MUXCY_L port map (
    DI => R1IN_4_ADD_1(9),
    CI => R1IN_4_ADD_2_0_CRY_8,
    S => R1IN_4_ADD_2_0_AXB_9,
    LO => R1IN_4_ADD_2_0_CRY_9);
R1IN_4_ADD_2_0_S_8: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_8,
    CI => R1IN_4_ADD_2_0_CRY_7,
    O => R1IN_4(25));
R1IN_4_ADD_2_0_CRY_8_Z8530: MUXCY_L port map (
    DI => R1IN_4_ADD_1(8),
    CI => R1IN_4_ADD_2_0_CRY_7,
    S => R1IN_4_ADD_2_0_AXB_8,
    LO => R1IN_4_ADD_2_0_CRY_8);
R1IN_4_ADD_2_0_S_7: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_7,
    CI => R1IN_4_ADD_2_0_CRY_6,
    O => R1IN_4(24));
R1IN_4_ADD_2_0_CRY_7_Z8532: MUXCY_L port map (
    DI => R1IN_4_ADD_1(7),
    CI => R1IN_4_ADD_2_0_CRY_6,
    S => R1IN_4_ADD_2_0_AXB_7,
    LO => R1IN_4_ADD_2_0_CRY_7);
R1IN_4_ADD_2_0_S_6: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_6,
    CI => R1IN_4_ADD_2_0_CRY_5,
    O => R1IN_4(23));
R1IN_4_ADD_2_0_CRY_6_Z8534: MUXCY_L port map (
    DI => R1IN_4_ADD_1(6),
    CI => R1IN_4_ADD_2_0_CRY_5,
    S => R1IN_4_ADD_2_0_AXB_6,
    LO => R1IN_4_ADD_2_0_CRY_6);
R1IN_4_ADD_2_0_S_5: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_5,
    CI => R1IN_4_ADD_2_0_CRY_4,
    O => R1IN_4(22));
R1IN_4_ADD_2_0_CRY_5_Z8536: MUXCY_L port map (
    DI => R1IN_4_ADD_1(5),
    CI => R1IN_4_ADD_2_0_CRY_4,
    S => R1IN_4_ADD_2_0_AXB_5,
    LO => R1IN_4_ADD_2_0_CRY_5);
R1IN_4_ADD_2_0_S_4: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_4,
    CI => R1IN_4_ADD_2_0_CRY_3,
    O => R1IN_4(21));
R1IN_4_ADD_2_0_CRY_4_Z8538: MUXCY_L port map (
    DI => R1IN_4_ADD_1(4),
    CI => R1IN_4_ADD_2_0_CRY_3,
    S => R1IN_4_ADD_2_0_AXB_4,
    LO => R1IN_4_ADD_2_0_CRY_4);
R1IN_4_ADD_2_0_S_3: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_3,
    CI => R1IN_4_ADD_2_0_CRY_2,
    O => R1IN_4(20));
R1IN_4_ADD_2_0_CRY_3_Z8540: MUXCY_L port map (
    DI => R1IN_4_ADD_1(3),
    CI => R1IN_4_ADD_2_0_CRY_2,
    S => R1IN_4_ADD_2_0_AXB_3,
    LO => R1IN_4_ADD_2_0_CRY_3);
R1IN_4_ADD_2_0_S_2: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_2,
    CI => R1IN_4_ADD_2_0_CRY_1,
    O => R1IN_4(19));
R1IN_4_ADD_2_0_CRY_2_Z8542: MUXCY_L port map (
    DI => R1IN_4_ADD_1(2),
    CI => R1IN_4_ADD_2_0_CRY_1,
    S => R1IN_4_ADD_2_0_AXB_2,
    LO => R1IN_4_ADD_2_0_CRY_2);
R1IN_4_ADD_2_0_S_1: XORCY port map (
    LI => R1IN_4_ADD_2_0_AXB_1,
    CI => R1IN_4_ADD_2_0_CRY_0,
    O => R1IN_4(18));
R1IN_4_ADD_2_0_CRY_1_Z8544: MUXCY_L port map (
    DI => R1IN_4_ADD_1(1),
    CI => R1IN_4_ADD_2_0_CRY_0,
    S => R1IN_4_ADD_2_0_AXB_1,
    LO => R1IN_4_ADD_2_0_CRY_1);
R1IN_4_ADD_2_0_CRY_0_Z8545: MUXCY_L port map (
    DI => R1IN_4_ADD_2_0,
    CI => NN_1,
    S => R1IN_4(17),
    LO => R1IN_4_ADD_2_0_CRY_0);
\R1IN_4_4_4[19:0]\: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 1,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => A(51),
  A(1) => A(52),
  A(2) => A(53),
  A(3) => A(54),
  A(4) => A(55),
  A(5) => A(56),
  A(6) => A(57),
  A(7) => A(58),
  A(8) => A(59),
  A(9) => A(60),
  A(10) => NN_1,
  A(11) => NN_1,
  A(12) => NN_1,
  A(13) => NN_1,
  A(14) => NN_1,
  A(15) => NN_1,
  A(16) => NN_1,
  A(17) => NN_1,
  B(0) => B(51),
  B(1) => B(52),
  B(2) => B(53),
  B(3) => B(54),
  B(4) => B(55),
  B(5) => B(56),
  B(6) => B(57),
  B(7) => B(58),
  B(8) => B(59),
  B(9) => B(60),
  B(10) => NN_1,
  B(11) => NN_1,
  B(12) => NN_1,
  B(13) => NN_1,
  B(14) => NN_1,
  B(15) => NN_1,
  B(16) => NN_1,
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => NN_1,
  PCIN(1) => NN_1,
  PCIN(2) => NN_1,
  PCIN(3) => NN_1,
  PCIN(4) => NN_1,
  PCIN(5) => NN_1,
  PCIN(6) => NN_1,
  PCIN(7) => NN_1,
  PCIN(8) => NN_1,
  PCIN(9) => NN_1,
  PCIN(10) => NN_1,
  PCIN(11) => NN_1,
  PCIN(12) => NN_1,
  PCIN(13) => NN_1,
  PCIN(14) => NN_1,
  PCIN(15) => NN_1,
  PCIN(16) => NN_1,
  PCIN(17) => NN_1,
  PCIN(18) => NN_1,
  PCIN(19) => NN_1,
  PCIN(20) => NN_1,
  PCIN(21) => NN_1,
  PCIN(22) => NN_1,
  PCIN(23) => NN_1,
  PCIN(24) => NN_1,
  PCIN(25) => NN_1,
  PCIN(26) => NN_1,
  PCIN(27) => NN_1,
  PCIN(28) => NN_1,
  PCIN(29) => NN_1,
  PCIN(30) => NN_1,
  PCIN(31) => NN_1,
  PCIN(32) => NN_1,
  PCIN(33) => NN_1,
  PCIN(34) => NN_1,
  PCIN(35) => NN_1,
  PCIN(36) => NN_1,
  PCIN(37) => NN_1,
  PCIN(38) => NN_1,
  PCIN(39) => NN_1,
  PCIN(40) => NN_1,
  PCIN(41) => NN_1,
  PCIN(42) => NN_1,
  PCIN(43) => NN_1,
  PCIN(44) => NN_1,
  PCIN(45) => NN_1,
  PCIN(46) => NN_1,
  PCIN(47) => NN_1,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_1,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => CLK,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => EN,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_4_4_4_BCOUT(0),
  BCOUT(1) => R1IN_4_4_4_BCOUT(1),
  BCOUT(2) => R1IN_4_4_4_BCOUT(2),
  BCOUT(3) => R1IN_4_4_4_BCOUT(3),
  BCOUT(4) => R1IN_4_4_4_BCOUT(4),
  BCOUT(5) => R1IN_4_4_4_BCOUT(5),
  BCOUT(6) => R1IN_4_4_4_BCOUT(6),
  BCOUT(7) => R1IN_4_4_4_BCOUT(7),
  BCOUT(8) => R1IN_4_4_4_BCOUT(8),
  BCOUT(9) => R1IN_4_4_4_BCOUT(9),
  BCOUT(10) => R1IN_4_4_4_BCOUT(10),
  BCOUT(11) => R1IN_4_4_4_BCOUT(11),
  BCOUT(12) => R1IN_4_4_4_BCOUT(12),
  BCOUT(13) => R1IN_4_4_4_BCOUT(13),
  BCOUT(14) => R1IN_4_4_4_BCOUT(14),
  BCOUT(15) => R1IN_4_4_4_BCOUT(15),
  BCOUT(16) => R1IN_4_4_4_BCOUT(16),
  BCOUT(17) => R1IN_4_4_4_BCOUT(17),
  P(0) => R1IN_4_4_4F(0),
  P(1) => R1IN_4_4_4F(1),
  P(2) => R1IN_4_4_4F(2),
  P(3) => R1IN_4_4_4F(3),
  P(4) => R1IN_4_4_4F(4),
  P(5) => R1IN_4_4_4F(5),
  P(6) => R1IN_4_4_4F(6),
  P(7) => R1IN_4_4_4F(7),
  P(8) => R1IN_4_4_4F(8),
  P(9) => R1IN_4_4_4F(9),
  P(10) => R1IN_4_4_4F(10),
  P(11) => R1IN_4_4_4F(11),
  P(12) => R1IN_4_4_4F(12),
  P(13) => R1IN_4_4_4F(13),
  P(14) => R1IN_4_4_4F(14),
  P(15) => R1IN_4_4_4F(15),
  P(16) => R1IN_4_4_4F(16),
  P(17) => R1IN_4_4_4F(17),
  P(18) => R1IN_4_4_4F(18),
  P(19) => R1IN_4_4_4F(19),
  P(20) => UC_250,
  P(21) => UC_251,
  P(22) => UC_252,
  P(23) => UC_253,
  P(24) => UC_254,
  P(25) => UC_255,
  P(26) => UC_256,
  P(27) => UC_257,
  P(28) => UC_258,
  P(29) => UC_259,
  P(30) => UC_260,
  P(31) => UC_261,
  P(32) => UC_262,
  P(33) => UC_263,
  P(34) => UC_264,
  P(35) => UC_265,
  P(36) => UC_266,
  P(37) => UC_267,
  P(38) => UC_268,
  P(39) => UC_269,
  P(40) => UC_270,
  P(41) => UC_271,
  P(42) => UC_272,
  P(43) => UC_273,
  P(44) => UC_274,
  P(45) => UC_275,
  P(46) => UC_276,
  P(47) => UC_277,
  PCOUT(0) => R1IN_4_4_4_PCOUT(0),
  PCOUT(1) => R1IN_4_4_4_PCOUT(1),
  PCOUT(2) => R1IN_4_4_4_PCOUT(2),
  PCOUT(3) => R1IN_4_4_4_PCOUT(3),
  PCOUT(4) => R1IN_4_4_4_PCOUT(4),
  PCOUT(5) => R1IN_4_4_4_PCOUT(5),
  PCOUT(6) => R1IN_4_4_4_PCOUT(6),
  PCOUT(7) => R1IN_4_4_4_PCOUT(7),
  PCOUT(8) => R1IN_4_4_4_PCOUT(8),
  PCOUT(9) => R1IN_4_4_4_PCOUT(9),
  PCOUT(10) => R1IN_4_4_4_PCOUT(10),
  PCOUT(11) => R1IN_4_4_4_PCOUT(11),
  PCOUT(12) => R1IN_4_4_4_PCOUT(12),
  PCOUT(13) => R1IN_4_4_4_PCOUT(13),
  PCOUT(14) => R1IN_4_4_4_PCOUT(14),
  PCOUT(15) => R1IN_4_4_4_PCOUT(15),
  PCOUT(16) => R1IN_4_4_4_PCOUT(16),
  PCOUT(17) => R1IN_4_4_4_PCOUT(17),
  PCOUT(18) => R1IN_4_4_4_PCOUT(18),
  PCOUT(19) => R1IN_4_4_4_PCOUT(19),
  PCOUT(20) => R1IN_4_4_4_PCOUT(20),
  PCOUT(21) => R1IN_4_4_4_PCOUT(21),
  PCOUT(22) => R1IN_4_4_4_PCOUT(22),
  PCOUT(23) => R1IN_4_4_4_PCOUT(23),
  PCOUT(24) => R1IN_4_4_4_PCOUT(24),
  PCOUT(25) => R1IN_4_4_4_PCOUT(25),
  PCOUT(26) => R1IN_4_4_4_PCOUT(26),
  PCOUT(27) => R1IN_4_4_4_PCOUT(27),
  PCOUT(28) => R1IN_4_4_4_PCOUT(28),
  PCOUT(29) => R1IN_4_4_4_PCOUT(29),
  PCOUT(30) => R1IN_4_4_4_PCOUT(30),
  PCOUT(31) => R1IN_4_4_4_PCOUT(31),
  PCOUT(32) => R1IN_4_4_4_PCOUT(32),
  PCOUT(33) => R1IN_4_4_4_PCOUT(33),
  PCOUT(34) => R1IN_4_4_4_PCOUT(34),
  PCOUT(35) => R1IN_4_4_4_PCOUT(35),
  PCOUT(36) => R1IN_4_4_4_PCOUT(36),
  PCOUT(37) => R1IN_4_4_4_PCOUT(37),
  PCOUT(38) => R1IN_4_4_4_PCOUT(38),
  PCOUT(39) => R1IN_4_4_4_PCOUT(39),
  PCOUT(40) => R1IN_4_4_4_PCOUT(40),
  PCOUT(41) => R1IN_4_4_4_PCOUT(41),
  PCOUT(42) => R1IN_4_4_4_PCOUT(42),
  PCOUT(43) => R1IN_4_4_4_PCOUT(43),
  PCOUT(44) => R1IN_4_4_4_PCOUT(44),
  PCOUT(45) => R1IN_4_4_4_PCOUT(45),
  PCOUT(46) => R1IN_4_4_4_PCOUT(46),
  PCOUT(47) => R1IN_4_4_4_PCOUT(47));
\R1IN_4_4_2[26:0]\: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 0,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => A(51),
  A(1) => A(52),
  A(2) => A(53),
  A(3) => A(54),
  A(4) => A(55),
  A(5) => A(56),
  A(6) => A(57),
  A(7) => A(58),
  A(8) => A(59),
  A(9) => A(60),
  A(10) => NN_1,
  A(11) => NN_1,
  A(12) => NN_1,
  A(13) => NN_1,
  A(14) => NN_1,
  A(15) => NN_1,
  A(16) => NN_1,
  A(17) => NN_1,
  B(0) => B(34),
  B(1) => B(35),
  B(2) => B(36),
  B(3) => B(37),
  B(4) => B(38),
  B(5) => B(39),
  B(6) => B(40),
  B(7) => B(41),
  B(8) => B(42),
  B(9) => B(43),
  B(10) => B(44),
  B(11) => B(45),
  B(12) => B(46),
  B(13) => B(47),
  B(14) => B(48),
  B(15) => B(49),
  B(16) => B(50),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => NN_1,
  PCIN(1) => NN_1,
  PCIN(2) => NN_1,
  PCIN(3) => NN_1,
  PCIN(4) => NN_1,
  PCIN(5) => NN_1,
  PCIN(6) => NN_1,
  PCIN(7) => NN_1,
  PCIN(8) => NN_1,
  PCIN(9) => NN_1,
  PCIN(10) => NN_1,
  PCIN(11) => NN_1,
  PCIN(12) => NN_1,
  PCIN(13) => NN_1,
  PCIN(14) => NN_1,
  PCIN(15) => NN_1,
  PCIN(16) => NN_1,
  PCIN(17) => NN_1,
  PCIN(18) => NN_1,
  PCIN(19) => NN_1,
  PCIN(20) => NN_1,
  PCIN(21) => NN_1,
  PCIN(22) => NN_1,
  PCIN(23) => NN_1,
  PCIN(24) => NN_1,
  PCIN(25) => NN_1,
  PCIN(26) => NN_1,
  PCIN(27) => NN_1,
  PCIN(28) => NN_1,
  PCIN(29) => NN_1,
  PCIN(30) => NN_1,
  PCIN(31) => NN_1,
  PCIN(32) => NN_1,
  PCIN(33) => NN_1,
  PCIN(34) => NN_1,
  PCIN(35) => NN_1,
  PCIN(36) => NN_1,
  PCIN(37) => NN_1,
  PCIN(38) => NN_1,
  PCIN(39) => NN_1,
  PCIN(40) => NN_1,
  PCIN(41) => NN_1,
  PCIN(42) => NN_1,
  PCIN(43) => NN_1,
  PCIN(44) => NN_1,
  PCIN(45) => NN_1,
  PCIN(46) => NN_1,
  PCIN(47) => NN_1,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_1,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => NN_1,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => NN_1,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_4_4_2_BCOUT(0),
  BCOUT(1) => R1IN_4_4_2_BCOUT(1),
  BCOUT(2) => R1IN_4_4_2_BCOUT(2),
  BCOUT(3) => R1IN_4_4_2_BCOUT(3),
  BCOUT(4) => R1IN_4_4_2_BCOUT(4),
  BCOUT(5) => R1IN_4_4_2_BCOUT(5),
  BCOUT(6) => R1IN_4_4_2_BCOUT(6),
  BCOUT(7) => R1IN_4_4_2_BCOUT(7),
  BCOUT(8) => R1IN_4_4_2_BCOUT(8),
  BCOUT(9) => R1IN_4_4_2_BCOUT(9),
  BCOUT(10) => R1IN_4_4_2_BCOUT(10),
  BCOUT(11) => R1IN_4_4_2_BCOUT(11),
  BCOUT(12) => R1IN_4_4_2_BCOUT(12),
  BCOUT(13) => R1IN_4_4_2_BCOUT(13),
  BCOUT(14) => R1IN_4_4_2_BCOUT(14),
  BCOUT(15) => R1IN_4_4_2_BCOUT(15),
  BCOUT(16) => R1IN_4_4_2_BCOUT(16),
  BCOUT(17) => R1IN_4_4_2_BCOUT(17),
  P(0) => R1IN_4_4_2(0),
  P(1) => R1IN_4_4_2(1),
  P(2) => R1IN_4_4_2(2),
  P(3) => R1IN_4_4_2(3),
  P(4) => R1IN_4_4_2(4),
  P(5) => R1IN_4_4_2(5),
  P(6) => R1IN_4_4_2(6),
  P(7) => R1IN_4_4_2(7),
  P(8) => R1IN_4_4_2(8),
  P(9) => R1IN_4_4_2(9),
  P(10) => R1IN_4_4_2(10),
  P(11) => R1IN_4_4_2(11),
  P(12) => R1IN_4_4_2(12),
  P(13) => R1IN_4_4_2(13),
  P(14) => R1IN_4_4_2(14),
  P(15) => R1IN_4_4_2(15),
  P(16) => R1IN_4_4_2(16),
  P(17) => R1IN_4_4_2(17),
  P(18) => R1IN_4_4_2(18),
  P(19) => R1IN_4_4_2(19),
  P(20) => R1IN_4_4_2(20),
  P(21) => R1IN_4_4_2(21),
  P(22) => R1IN_4_4_2(22),
  P(23) => R1IN_4_4_2(23),
  P(24) => R1IN_4_4_2(24),
  P(25) => R1IN_4_4_2(25),
  P(26) => R1IN_4_4_2(26),
  P(27) => UC_229,
  P(28) => UC_230,
  P(29) => UC_231,
  P(30) => UC_232,
  P(31) => UC_233,
  P(32) => UC_234,
  P(33) => UC_235,
  P(34) => UC_236,
  P(35) => UC_237,
  P(36) => UC_238,
  P(37) => UC_239,
  P(38) => UC_240,
  P(39) => UC_241,
  P(40) => UC_242,
  P(41) => UC_243,
  P(42) => UC_244,
  P(43) => UC_245,
  P(44) => UC_246,
  P(45) => UC_247,
  P(46) => UC_248,
  P(47) => UC_249,
  PCOUT(0) => R1IN_4_4_2_0(0),
  PCOUT(1) => R1IN_4_4_2_0(1),
  PCOUT(2) => R1IN_4_4_2_0(2),
  PCOUT(3) => R1IN_4_4_2_0(3),
  PCOUT(4) => R1IN_4_4_2_0(4),
  PCOUT(5) => R1IN_4_4_2_0(5),
  PCOUT(6) => R1IN_4_4_2_0(6),
  PCOUT(7) => R1IN_4_4_2_0(7),
  PCOUT(8) => R1IN_4_4_2_0(8),
  PCOUT(9) => R1IN_4_4_2_0(9),
  PCOUT(10) => R1IN_4_4_2_0(10),
  PCOUT(11) => R1IN_4_4_2_0(11),
  PCOUT(12) => R1IN_4_4_2_0(12),
  PCOUT(13) => R1IN_4_4_2_0(13),
  PCOUT(14) => R1IN_4_4_2_0(14),
  PCOUT(15) => R1IN_4_4_2_0(15),
  PCOUT(16) => R1IN_4_4_2_0(16),
  PCOUT(17) => R1IN_4_4_2_0(17),
  PCOUT(18) => R1IN_4_4_2_0(18),
  PCOUT(19) => R1IN_4_4_2_0(19),
  PCOUT(20) => R1IN_4_4_2_0(20),
  PCOUT(21) => R1IN_4_4_2_0(21),
  PCOUT(22) => R1IN_4_4_2_0(22),
  PCOUT(23) => R1IN_4_4_2_0(23),
  PCOUT(24) => R1IN_4_4_2_0(24),
  PCOUT(25) => R1IN_4_4_2_0(25),
  PCOUT(26) => R1IN_4_4_2_0(26),
  PCOUT(27) => UC_229_0,
  PCOUT(28) => UC_230_0,
  PCOUT(29) => UC_231_0,
  PCOUT(30) => UC_232_0,
  PCOUT(31) => UC_233_0,
  PCOUT(32) => UC_234_0,
  PCOUT(33) => UC_235_0,
  PCOUT(34) => UC_236_0,
  PCOUT(35) => UC_237_0,
  PCOUT(36) => UC_238_0,
  PCOUT(37) => UC_239_0,
  PCOUT(38) => UC_240_0,
  PCOUT(39) => UC_241_0,
  PCOUT(40) => UC_242_0,
  PCOUT(41) => UC_243_0,
  PCOUT(42) => UC_244_0,
  PCOUT(43) => UC_245_0,
  PCOUT(44) => UC_246_0,
  PCOUT(45) => UC_247_0,
  PCOUT(46) => UC_248_0,
  PCOUT(47) => UC_249_0);
\R1IN_4_4_1[33:0]\: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 1,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => A(34),
  A(1) => A(35),
  A(2) => A(36),
  A(3) => A(37),
  A(4) => A(38),
  A(5) => A(39),
  A(6) => A(40),
  A(7) => A(41),
  A(8) => A(42),
  A(9) => A(43),
  A(10) => A(44),
  A(11) => A(45),
  A(12) => A(46),
  A(13) => A(47),
  A(14) => A(48),
  A(15) => A(49),
  A(16) => A(50),
  A(17) => NN_1,
  B(0) => B(34),
  B(1) => B(35),
  B(2) => B(36),
  B(3) => B(37),
  B(4) => B(38),
  B(5) => B(39),
  B(6) => B(40),
  B(7) => B(41),
  B(8) => B(42),
  B(9) => B(43),
  B(10) => B(44),
  B(11) => B(45),
  B(12) => B(46),
  B(13) => B(47),
  B(14) => B(48),
  B(15) => B(49),
  B(16) => B(50),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => NN_1,
  PCIN(1) => NN_1,
  PCIN(2) => NN_1,
  PCIN(3) => NN_1,
  PCIN(4) => NN_1,
  PCIN(5) => NN_1,
  PCIN(6) => NN_1,
  PCIN(7) => NN_1,
  PCIN(8) => NN_1,
  PCIN(9) => NN_1,
  PCIN(10) => NN_1,
  PCIN(11) => NN_1,
  PCIN(12) => NN_1,
  PCIN(13) => NN_1,
  PCIN(14) => NN_1,
  PCIN(15) => NN_1,
  PCIN(16) => NN_1,
  PCIN(17) => NN_1,
  PCIN(18) => NN_1,
  PCIN(19) => NN_1,
  PCIN(20) => NN_1,
  PCIN(21) => NN_1,
  PCIN(22) => NN_1,
  PCIN(23) => NN_1,
  PCIN(24) => NN_1,
  PCIN(25) => NN_1,
  PCIN(26) => NN_1,
  PCIN(27) => NN_1,
  PCIN(28) => NN_1,
  PCIN(29) => NN_1,
  PCIN(30) => NN_1,
  PCIN(31) => NN_1,
  PCIN(32) => NN_1,
  PCIN(33) => NN_1,
  PCIN(34) => NN_1,
  PCIN(35) => NN_1,
  PCIN(36) => NN_1,
  PCIN(37) => NN_1,
  PCIN(38) => NN_1,
  PCIN(39) => NN_1,
  PCIN(40) => NN_1,
  PCIN(41) => NN_1,
  PCIN(42) => NN_1,
  PCIN(43) => NN_1,
  PCIN(44) => NN_1,
  PCIN(45) => NN_1,
  PCIN(46) => NN_1,
  PCIN(47) => NN_1,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_1,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => CLK,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => EN,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_4_4_1_BCOUT(0),
  BCOUT(1) => R1IN_4_4_1_BCOUT(1),
  BCOUT(2) => R1IN_4_4_1_BCOUT(2),
  BCOUT(3) => R1IN_4_4_1_BCOUT(3),
  BCOUT(4) => R1IN_4_4_1_BCOUT(4),
  BCOUT(5) => R1IN_4_4_1_BCOUT(5),
  BCOUT(6) => R1IN_4_4_1_BCOUT(6),
  BCOUT(7) => R1IN_4_4_1_BCOUT(7),
  BCOUT(8) => R1IN_4_4_1_BCOUT(8),
  BCOUT(9) => R1IN_4_4_1_BCOUT(9),
  BCOUT(10) => R1IN_4_4_1_BCOUT(10),
  BCOUT(11) => R1IN_4_4_1_BCOUT(11),
  BCOUT(12) => R1IN_4_4_1_BCOUT(12),
  BCOUT(13) => R1IN_4_4_1_BCOUT(13),
  BCOUT(14) => R1IN_4_4_1_BCOUT(14),
  BCOUT(15) => R1IN_4_4_1_BCOUT(15),
  BCOUT(16) => R1IN_4_4_1_BCOUT(16),
  BCOUT(17) => R1IN_4_4_1_BCOUT(17),
  P(0) => R1IN_4_4F(0),
  P(1) => R1IN_4_4F(1),
  P(2) => R1IN_4_4F(2),
  P(3) => R1IN_4_4F(3),
  P(4) => R1IN_4_4F(4),
  P(5) => R1IN_4_4F(5),
  P(6) => R1IN_4_4F(6),
  P(7) => R1IN_4_4F(7),
  P(8) => R1IN_4_4F(8),
  P(9) => R1IN_4_4F(9),
  P(10) => R1IN_4_4F(10),
  P(11) => R1IN_4_4F(11),
  P(12) => R1IN_4_4F(12),
  P(13) => R1IN_4_4F(13),
  P(14) => R1IN_4_4F(14),
  P(15) => R1IN_4_4F(15),
  P(16) => R1IN_4_4F(16),
  P(17) => R1IN_4_4_ADD_2,
  P(18) => R1IN_4_4_1F(18),
  P(19) => R1IN_4_4_1F(19),
  P(20) => R1IN_4_4_1F(20),
  P(21) => R1IN_4_4_1F(21),
  P(22) => R1IN_4_4_1F(22),
  P(23) => R1IN_4_4_1F(23),
  P(24) => R1IN_4_4_1F(24),
  P(25) => R1IN_4_4_1F(25),
  P(26) => R1IN_4_4_1F(26),
  P(27) => R1IN_4_4_1F(27),
  P(28) => R1IN_4_4_1F(28),
  P(29) => R1IN_4_4_1F(29),
  P(30) => R1IN_4_4_1F(30),
  P(31) => R1IN_4_4_1F(31),
  P(32) => R1IN_4_4_1F(32),
  P(33) => R1IN_4_4_1F(33),
  P(34) => UC_215,
  P(35) => UC_216,
  P(36) => UC_217,
  P(37) => UC_218,
  P(38) => UC_219,
  P(39) => UC_220,
  P(40) => UC_221,
  P(41) => UC_222,
  P(42) => UC_223,
  P(43) => UC_224,
  P(44) => UC_225,
  P(45) => UC_226,
  P(46) => UC_227,
  P(47) => UC_228,
  PCOUT(0) => R1IN_4_4_1_PCOUT(0),
  PCOUT(1) => R1IN_4_4_1_PCOUT(1),
  PCOUT(2) => R1IN_4_4_1_PCOUT(2),
  PCOUT(3) => R1IN_4_4_1_PCOUT(3),
  PCOUT(4) => R1IN_4_4_1_PCOUT(4),
  PCOUT(5) => R1IN_4_4_1_PCOUT(5),
  PCOUT(6) => R1IN_4_4_1_PCOUT(6),
  PCOUT(7) => R1IN_4_4_1_PCOUT(7),
  PCOUT(8) => R1IN_4_4_1_PCOUT(8),
  PCOUT(9) => R1IN_4_4_1_PCOUT(9),
  PCOUT(10) => R1IN_4_4_1_PCOUT(10),
  PCOUT(11) => R1IN_4_4_1_PCOUT(11),
  PCOUT(12) => R1IN_4_4_1_PCOUT(12),
  PCOUT(13) => R1IN_4_4_1_PCOUT(13),
  PCOUT(14) => R1IN_4_4_1_PCOUT(14),
  PCOUT(15) => R1IN_4_4_1_PCOUT(15),
  PCOUT(16) => R1IN_4_4_1_PCOUT(16),
  PCOUT(17) => R1IN_4_4_1_PCOUT(17),
  PCOUT(18) => R1IN_4_4_1_PCOUT(18),
  PCOUT(19) => R1IN_4_4_1_PCOUT(19),
  PCOUT(20) => R1IN_4_4_1_PCOUT(20),
  PCOUT(21) => R1IN_4_4_1_PCOUT(21),
  PCOUT(22) => R1IN_4_4_1_PCOUT(22),
  PCOUT(23) => R1IN_4_4_1_PCOUT(23),
  PCOUT(24) => R1IN_4_4_1_PCOUT(24),
  PCOUT(25) => R1IN_4_4_1_PCOUT(25),
  PCOUT(26) => R1IN_4_4_1_PCOUT(26),
  PCOUT(27) => R1IN_4_4_1_PCOUT(27),
  PCOUT(28) => R1IN_4_4_1_PCOUT(28),
  PCOUT(29) => R1IN_4_4_1_PCOUT(29),
  PCOUT(30) => R1IN_4_4_1_PCOUT(30),
  PCOUT(31) => R1IN_4_4_1_PCOUT(31),
  PCOUT(32) => R1IN_4_4_1_PCOUT(32),
  PCOUT(33) => R1IN_4_4_1_PCOUT(33),
  PCOUT(34) => R1IN_4_4_1_PCOUT(34),
  PCOUT(35) => R1IN_4_4_1_PCOUT(35),
  PCOUT(36) => R1IN_4_4_1_PCOUT(36),
  PCOUT(37) => R1IN_4_4_1_PCOUT(37),
  PCOUT(38) => R1IN_4_4_1_PCOUT(38),
  PCOUT(39) => R1IN_4_4_1_PCOUT(39),
  PCOUT(40) => R1IN_4_4_1_PCOUT(40),
  PCOUT(41) => R1IN_4_4_1_PCOUT(41),
  PCOUT(42) => R1IN_4_4_1_PCOUT(42),
  PCOUT(43) => R1IN_4_4_1_PCOUT(43),
  PCOUT(44) => R1IN_4_4_1_PCOUT(44),
  PCOUT(45) => R1IN_4_4_1_PCOUT(45),
  PCOUT(46) => R1IN_4_4_1_PCOUT(46),
  PCOUT(47) => R1IN_4_4_1_PCOUT(47));
\R1IN_4_1[33:0]\: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 1,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => A(17),
  A(1) => A(18),
  A(2) => A(19),
  A(3) => A(20),
  A(4) => A(21),
  A(5) => A(22),
  A(6) => A(23),
  A(7) => A(24),
  A(8) => A(25),
  A(9) => A(26),
  A(10) => A(27),
  A(11) => A(28),
  A(12) => A(29),
  A(13) => A(30),
  A(14) => A(31),
  A(15) => A(32),
  A(16) => A(33),
  A(17) => NN_1,
  B(0) => B(17),
  B(1) => B(18),
  B(2) => B(19),
  B(3) => B(20),
  B(4) => B(21),
  B(5) => B(22),
  B(6) => B(23),
  B(7) => B(24),
  B(8) => B(25),
  B(9) => B(26),
  B(10) => B(27),
  B(11) => B(28),
  B(12) => B(29),
  B(13) => B(30),
  B(14) => B(31),
  B(15) => B(32),
  B(16) => B(33),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => NN_1,
  PCIN(1) => NN_1,
  PCIN(2) => NN_1,
  PCIN(3) => NN_1,
  PCIN(4) => NN_1,
  PCIN(5) => NN_1,
  PCIN(6) => NN_1,
  PCIN(7) => NN_1,
  PCIN(8) => NN_1,
  PCIN(9) => NN_1,
  PCIN(10) => NN_1,
  PCIN(11) => NN_1,
  PCIN(12) => NN_1,
  PCIN(13) => NN_1,
  PCIN(14) => NN_1,
  PCIN(15) => NN_1,
  PCIN(16) => NN_1,
  PCIN(17) => NN_1,
  PCIN(18) => NN_1,
  PCIN(19) => NN_1,
  PCIN(20) => NN_1,
  PCIN(21) => NN_1,
  PCIN(22) => NN_1,
  PCIN(23) => NN_1,
  PCIN(24) => NN_1,
  PCIN(25) => NN_1,
  PCIN(26) => NN_1,
  PCIN(27) => NN_1,
  PCIN(28) => NN_1,
  PCIN(29) => NN_1,
  PCIN(30) => NN_1,
  PCIN(31) => NN_1,
  PCIN(32) => NN_1,
  PCIN(33) => NN_1,
  PCIN(34) => NN_1,
  PCIN(35) => NN_1,
  PCIN(36) => NN_1,
  PCIN(37) => NN_1,
  PCIN(38) => NN_1,
  PCIN(39) => NN_1,
  PCIN(40) => NN_1,
  PCIN(41) => NN_1,
  PCIN(42) => NN_1,
  PCIN(43) => NN_1,
  PCIN(44) => NN_1,
  PCIN(45) => NN_1,
  PCIN(46) => NN_1,
  PCIN(47) => NN_1,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_1,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => CLK,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => EN,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_4_1_BCOUT(0),
  BCOUT(1) => R1IN_4_1_BCOUT(1),
  BCOUT(2) => R1IN_4_1_BCOUT(2),
  BCOUT(3) => R1IN_4_1_BCOUT(3),
  BCOUT(4) => R1IN_4_1_BCOUT(4),
  BCOUT(5) => R1IN_4_1_BCOUT(5),
  BCOUT(6) => R1IN_4_1_BCOUT(6),
  BCOUT(7) => R1IN_4_1_BCOUT(7),
  BCOUT(8) => R1IN_4_1_BCOUT(8),
  BCOUT(9) => R1IN_4_1_BCOUT(9),
  BCOUT(10) => R1IN_4_1_BCOUT(10),
  BCOUT(11) => R1IN_4_1_BCOUT(11),
  BCOUT(12) => R1IN_4_1_BCOUT(12),
  BCOUT(13) => R1IN_4_1_BCOUT(13),
  BCOUT(14) => R1IN_4_1_BCOUT(14),
  BCOUT(15) => R1IN_4_1_BCOUT(15),
  BCOUT(16) => R1IN_4_1_BCOUT(16),
  BCOUT(17) => R1IN_4_1_BCOUT(17),
  P(0) => R1IN_4F(0),
  P(1) => R1IN_4F(1),
  P(2) => R1IN_4F(2),
  P(3) => R1IN_4F(3),
  P(4) => R1IN_4F(4),
  P(5) => R1IN_4F(5),
  P(6) => R1IN_4F(6),
  P(7) => R1IN_4F(7),
  P(8) => R1IN_4F(8),
  P(9) => R1IN_4F(9),
  P(10) => R1IN_4F(10),
  P(11) => R1IN_4F(11),
  P(12) => R1IN_4F(12),
  P(13) => R1IN_4F(13),
  P(14) => R1IN_4F(14),
  P(15) => R1IN_4F(15),
  P(16) => R1IN_4F(16),
  P(17) => R1IN_4_1F(17),
  P(18) => R1IN_4_1F(18),
  P(19) => R1IN_4_1F(19),
  P(20) => R1IN_4_1F(20),
  P(21) => R1IN_4_1F(21),
  P(22) => R1IN_4_1F(22),
  P(23) => R1IN_4_1F(23),
  P(24) => R1IN_4_1F(24),
  P(25) => R1IN_4_1F(25),
  P(26) => R1IN_4_1F(26),
  P(27) => R1IN_4_1F(27),
  P(28) => R1IN_4_1F(28),
  P(29) => R1IN_4_1F(29),
  P(30) => R1IN_4_1F(30),
  P(31) => R1IN_4_1F(31),
  P(32) => R1IN_4_1F(32),
  P(33) => R1IN_4_1F(33),
  P(34) => UC_201,
  P(35) => UC_202,
  P(36) => UC_203,
  P(37) => UC_204,
  P(38) => UC_205,
  P(39) => UC_206,
  P(40) => UC_207,
  P(41) => UC_208,
  P(42) => UC_209,
  P(43) => UC_210,
  P(44) => UC_211,
  P(45) => UC_212,
  P(46) => UC_213,
  P(47) => UC_214,
  PCOUT(0) => R1IN_4_1_PCOUT(0),
  PCOUT(1) => R1IN_4_1_PCOUT(1),
  PCOUT(2) => R1IN_4_1_PCOUT(2),
  PCOUT(3) => R1IN_4_1_PCOUT(3),
  PCOUT(4) => R1IN_4_1_PCOUT(4),
  PCOUT(5) => R1IN_4_1_PCOUT(5),
  PCOUT(6) => R1IN_4_1_PCOUT(6),
  PCOUT(7) => R1IN_4_1_PCOUT(7),
  PCOUT(8) => R1IN_4_1_PCOUT(8),
  PCOUT(9) => R1IN_4_1_PCOUT(9),
  PCOUT(10) => R1IN_4_1_PCOUT(10),
  PCOUT(11) => R1IN_4_1_PCOUT(11),
  PCOUT(12) => R1IN_4_1_PCOUT(12),
  PCOUT(13) => R1IN_4_1_PCOUT(13),
  PCOUT(14) => R1IN_4_1_PCOUT(14),
  PCOUT(15) => R1IN_4_1_PCOUT(15),
  PCOUT(16) => R1IN_4_1_PCOUT(16),
  PCOUT(17) => R1IN_4_1_PCOUT(17),
  PCOUT(18) => R1IN_4_1_PCOUT(18),
  PCOUT(19) => R1IN_4_1_PCOUT(19),
  PCOUT(20) => R1IN_4_1_PCOUT(20),
  PCOUT(21) => R1IN_4_1_PCOUT(21),
  PCOUT(22) => R1IN_4_1_PCOUT(22),
  PCOUT(23) => R1IN_4_1_PCOUT(23),
  PCOUT(24) => R1IN_4_1_PCOUT(24),
  PCOUT(25) => R1IN_4_1_PCOUT(25),
  PCOUT(26) => R1IN_4_1_PCOUT(26),
  PCOUT(27) => R1IN_4_1_PCOUT(27),
  PCOUT(28) => R1IN_4_1_PCOUT(28),
  PCOUT(29) => R1IN_4_1_PCOUT(29),
  PCOUT(30) => R1IN_4_1_PCOUT(30),
  PCOUT(31) => R1IN_4_1_PCOUT(31),
  PCOUT(32) => R1IN_4_1_PCOUT(32),
  PCOUT(33) => R1IN_4_1_PCOUT(33),
  PCOUT(34) => R1IN_4_1_PCOUT(34),
  PCOUT(35) => R1IN_4_1_PCOUT(35),
  PCOUT(36) => R1IN_4_1_PCOUT(36),
  PCOUT(37) => R1IN_4_1_PCOUT(37),
  PCOUT(38) => R1IN_4_1_PCOUT(38),
  PCOUT(39) => R1IN_4_1_PCOUT(39),
  PCOUT(40) => R1IN_4_1_PCOUT(40),
  PCOUT(41) => R1IN_4_1_PCOUT(41),
  PCOUT(42) => R1IN_4_1_PCOUT(42),
  PCOUT(43) => R1IN_4_1_PCOUT(43),
  PCOUT(44) => R1IN_4_1_PCOUT(44),
  PCOUT(45) => R1IN_4_1_PCOUT(45),
  PCOUT(46) => R1IN_4_1_PCOUT(46),
  PCOUT(47) => R1IN_4_1_PCOUT(47));
\R1IN_3_1[33:0]\: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 0,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => B(17),
  A(1) => B(18),
  A(2) => B(19),
  A(3) => B(20),
  A(4) => B(21),
  A(5) => B(22),
  A(6) => B(23),
  A(7) => B(24),
  A(8) => B(25),
  A(9) => B(26),
  A(10) => B(27),
  A(11) => B(28),
  A(12) => B(29),
  A(13) => B(30),
  A(14) => B(31),
  A(15) => B(32),
  A(16) => B(33),
  A(17) => NN_1,
  B(0) => A(0),
  B(1) => A(1),
  B(2) => A(2),
  B(3) => A(3),
  B(4) => A(4),
  B(5) => A(5),
  B(6) => A(6),
  B(7) => A(7),
  B(8) => A(8),
  B(9) => A(9),
  B(10) => A(10),
  B(11) => A(11),
  B(12) => A(12),
  B(13) => A(13),
  B(14) => A(14),
  B(15) => A(15),
  B(16) => A(16),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => NN_1,
  PCIN(1) => NN_1,
  PCIN(2) => NN_1,
  PCIN(3) => NN_1,
  PCIN(4) => NN_1,
  PCIN(5) => NN_1,
  PCIN(6) => NN_1,
  PCIN(7) => NN_1,
  PCIN(8) => NN_1,
  PCIN(9) => NN_1,
  PCIN(10) => NN_1,
  PCIN(11) => NN_1,
  PCIN(12) => NN_1,
  PCIN(13) => NN_1,
  PCIN(14) => NN_1,
  PCIN(15) => NN_1,
  PCIN(16) => NN_1,
  PCIN(17) => NN_1,
  PCIN(18) => NN_1,
  PCIN(19) => NN_1,
  PCIN(20) => NN_1,
  PCIN(21) => NN_1,
  PCIN(22) => NN_1,
  PCIN(23) => NN_1,
  PCIN(24) => NN_1,
  PCIN(25) => NN_1,
  PCIN(26) => NN_1,
  PCIN(27) => NN_1,
  PCIN(28) => NN_1,
  PCIN(29) => NN_1,
  PCIN(30) => NN_1,
  PCIN(31) => NN_1,
  PCIN(32) => NN_1,
  PCIN(33) => NN_1,
  PCIN(34) => NN_1,
  PCIN(35) => NN_1,
  PCIN(36) => NN_1,
  PCIN(37) => NN_1,
  PCIN(38) => NN_1,
  PCIN(39) => NN_1,
  PCIN(40) => NN_1,
  PCIN(41) => NN_1,
  PCIN(42) => NN_1,
  PCIN(43) => NN_1,
  PCIN(44) => NN_1,
  PCIN(45) => NN_1,
  PCIN(46) => NN_1,
  PCIN(47) => NN_1,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_1,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => CLK,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => NN_1,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_3_1_BCOUT(0),
  BCOUT(1) => R1IN_3_1_BCOUT(1),
  BCOUT(2) => R1IN_3_1_BCOUT(2),
  BCOUT(3) => R1IN_3_1_BCOUT(3),
  BCOUT(4) => R1IN_3_1_BCOUT(4),
  BCOUT(5) => R1IN_3_1_BCOUT(5),
  BCOUT(6) => R1IN_3_1_BCOUT(6),
  BCOUT(7) => R1IN_3_1_BCOUT(7),
  BCOUT(8) => R1IN_3_1_BCOUT(8),
  BCOUT(9) => R1IN_3_1_BCOUT(9),
  BCOUT(10) => R1IN_3_1_BCOUT(10),
  BCOUT(11) => R1IN_3_1_BCOUT(11),
  BCOUT(12) => R1IN_3_1_BCOUT(12),
  BCOUT(13) => R1IN_3_1_BCOUT(13),
  BCOUT(14) => R1IN_3_1_BCOUT(14),
  BCOUT(15) => R1IN_3_1_BCOUT(15),
  BCOUT(16) => R1IN_3_1_BCOUT(16),
  BCOUT(17) => R1IN_3_1_BCOUT(17),
  P(0) => R1IN_3F_0(0),
  P(1) => R1IN_3F_0(1),
  P(2) => R1IN_3F_0(2),
  P(3) => R1IN_3F_0(3),
  P(4) => R1IN_3F_0(4),
  P(5) => R1IN_3F_0(5),
  P(6) => R1IN_3F_0(6),
  P(7) => R1IN_3F_0(7),
  P(8) => R1IN_3F_0(8),
  P(9) => R1IN_3F_0(9),
  P(10) => R1IN_3F_0(10),
  P(11) => R1IN_3F_0(11),
  P(12) => R1IN_3F_0(12),
  P(13) => R1IN_3F_0(13),
  P(14) => R1IN_3F_0(14),
  P(15) => R1IN_3F_0(15),
  P(16) => R1IN_3F_0(16),
  P(17) => R1IN_3_1F_0(17),
  P(18) => R1IN_3_1F_0(18),
  P(19) => R1IN_3_1F_0(19),
  P(20) => R1IN_3_1F_0(20),
  P(21) => R1IN_3_1F_0(21),
  P(22) => R1IN_3_1F_0(22),
  P(23) => R1IN_3_1F_0(23),
  P(24) => R1IN_3_1F_0(24),
  P(25) => R1IN_3_1F_0(25),
  P(26) => R1IN_3_1F_0(26),
  P(27) => R1IN_3_1F_0(27),
  P(28) => R1IN_3_1F_0(28),
  P(29) => R1IN_3_1F_0(29),
  P(30) => R1IN_3_1F_0(30),
  P(31) => R1IN_3_1F_0(31),
  P(32) => R1IN_3_1F_0(32),
  P(33) => R1IN_3_1F_0(33),
  P(34) => UC_187_0,
  P(35) => UC_188_0,
  P(36) => UC_189_0,
  P(37) => UC_190_0,
  P(38) => UC_191_0,
  P(39) => UC_192_0,
  P(40) => UC_193_0,
  P(41) => UC_194_0,
  P(42) => UC_195_0,
  P(43) => UC_196_0,
  P(44) => UC_197_0,
  P(45) => UC_198_0,
  P(46) => UC_199_0,
  P(47) => UC_200_0,
  PCOUT(0) => R1IN_3_1_PCOUT(0),
  PCOUT(1) => R1IN_3_1_PCOUT(1),
  PCOUT(2) => R1IN_3_1_PCOUT(2),
  PCOUT(3) => R1IN_3_1_PCOUT(3),
  PCOUT(4) => R1IN_3_1_PCOUT(4),
  PCOUT(5) => R1IN_3_1_PCOUT(5),
  PCOUT(6) => R1IN_3_1_PCOUT(6),
  PCOUT(7) => R1IN_3_1_PCOUT(7),
  PCOUT(8) => R1IN_3_1_PCOUT(8),
  PCOUT(9) => R1IN_3_1_PCOUT(9),
  PCOUT(10) => R1IN_3_1_PCOUT(10),
  PCOUT(11) => R1IN_3_1_PCOUT(11),
  PCOUT(12) => R1IN_3_1_PCOUT(12),
  PCOUT(13) => R1IN_3_1_PCOUT(13),
  PCOUT(14) => R1IN_3_1_PCOUT(14),
  PCOUT(15) => R1IN_3_1_PCOUT(15),
  PCOUT(16) => R1IN_3_1_PCOUT(16),
  PCOUT(17) => R1IN_3_1_PCOUT(17),
  PCOUT(18) => R1IN_3_1_PCOUT(18),
  PCOUT(19) => R1IN_3_1_PCOUT(19),
  PCOUT(20) => R1IN_3_1_PCOUT(20),
  PCOUT(21) => R1IN_3_1_PCOUT(21),
  PCOUT(22) => R1IN_3_1_PCOUT(22),
  PCOUT(23) => R1IN_3_1_PCOUT(23),
  PCOUT(24) => R1IN_3_1_PCOUT(24),
  PCOUT(25) => R1IN_3_1_PCOUT(25),
  PCOUT(26) => R1IN_3_1_PCOUT(26),
  PCOUT(27) => R1IN_3_1_PCOUT(27),
  PCOUT(28) => R1IN_3_1_PCOUT(28),
  PCOUT(29) => R1IN_3_1_PCOUT(29),
  PCOUT(30) => R1IN_3_1_PCOUT(30),
  PCOUT(31) => R1IN_3_1_PCOUT(31),
  PCOUT(32) => R1IN_3_1_PCOUT(32),
  PCOUT(33) => R1IN_3_1_PCOUT(33),
  PCOUT(34) => R1IN_3_1_PCOUT(34),
  PCOUT(35) => R1IN_3_1_PCOUT(35),
  PCOUT(36) => R1IN_3_1_PCOUT(36),
  PCOUT(37) => R1IN_3_1_PCOUT(37),
  PCOUT(38) => R1IN_3_1_PCOUT(38),
  PCOUT(39) => R1IN_3_1_PCOUT(39),
  PCOUT(40) => R1IN_3_1_PCOUT(40),
  PCOUT(41) => R1IN_3_1_PCOUT(41),
  PCOUT(42) => R1IN_3_1_PCOUT(42),
  PCOUT(43) => R1IN_3_1_PCOUT(43),
  PCOUT(44) => R1IN_3_1_PCOUT(44),
  PCOUT(45) => R1IN_3_1_PCOUT(45),
  PCOUT(46) => R1IN_3_1_PCOUT(46),
  PCOUT(47) => R1IN_3_1_PCOUT(47));
\R1IN_2_1[33:0]\: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 0,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => A(17),
  A(1) => A(18),
  A(2) => A(19),
  A(3) => A(20),
  A(4) => A(21),
  A(5) => A(22),
  A(6) => A(23),
  A(7) => A(24),
  A(8) => A(25),
  A(9) => A(26),
  A(10) => A(27),
  A(11) => A(28),
  A(12) => A(29),
  A(13) => A(30),
  A(14) => A(31),
  A(15) => A(32),
  A(16) => A(33),
  A(17) => NN_1,
  B(0) => B(0),
  B(1) => B(1),
  B(2) => B(2),
  B(3) => B(3),
  B(4) => B(4),
  B(5) => B(5),
  B(6) => B(6),
  B(7) => B(7),
  B(8) => B(8),
  B(9) => B(9),
  B(10) => B(10),
  B(11) => B(11),
  B(12) => B(12),
  B(13) => B(13),
  B(14) => B(14),
  B(15) => B(15),
  B(16) => B(16),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => NN_1,
  PCIN(1) => NN_1,
  PCIN(2) => NN_1,
  PCIN(3) => NN_1,
  PCIN(4) => NN_1,
  PCIN(5) => NN_1,
  PCIN(6) => NN_1,
  PCIN(7) => NN_1,
  PCIN(8) => NN_1,
  PCIN(9) => NN_1,
  PCIN(10) => NN_1,
  PCIN(11) => NN_1,
  PCIN(12) => NN_1,
  PCIN(13) => NN_1,
  PCIN(14) => NN_1,
  PCIN(15) => NN_1,
  PCIN(16) => NN_1,
  PCIN(17) => NN_1,
  PCIN(18) => NN_1,
  PCIN(19) => NN_1,
  PCIN(20) => NN_1,
  PCIN(21) => NN_1,
  PCIN(22) => NN_1,
  PCIN(23) => NN_1,
  PCIN(24) => NN_1,
  PCIN(25) => NN_1,
  PCIN(26) => NN_1,
  PCIN(27) => NN_1,
  PCIN(28) => NN_1,
  PCIN(29) => NN_1,
  PCIN(30) => NN_1,
  PCIN(31) => NN_1,
  PCIN(32) => NN_1,
  PCIN(33) => NN_1,
  PCIN(34) => NN_1,
  PCIN(35) => NN_1,
  PCIN(36) => NN_1,
  PCIN(37) => NN_1,
  PCIN(38) => NN_1,
  PCIN(39) => NN_1,
  PCIN(40) => NN_1,
  PCIN(41) => NN_1,
  PCIN(42) => NN_1,
  PCIN(43) => NN_1,
  PCIN(44) => NN_1,
  PCIN(45) => NN_1,
  PCIN(46) => NN_1,
  PCIN(47) => NN_1,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_1,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => CLK,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => NN_1,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_2_1_BCOUT(0),
  BCOUT(1) => R1IN_2_1_BCOUT(1),
  BCOUT(2) => R1IN_2_1_BCOUT(2),
  BCOUT(3) => R1IN_2_1_BCOUT(3),
  BCOUT(4) => R1IN_2_1_BCOUT(4),
  BCOUT(5) => R1IN_2_1_BCOUT(5),
  BCOUT(6) => R1IN_2_1_BCOUT(6),
  BCOUT(7) => R1IN_2_1_BCOUT(7),
  BCOUT(8) => R1IN_2_1_BCOUT(8),
  BCOUT(9) => R1IN_2_1_BCOUT(9),
  BCOUT(10) => R1IN_2_1_BCOUT(10),
  BCOUT(11) => R1IN_2_1_BCOUT(11),
  BCOUT(12) => R1IN_2_1_BCOUT(12),
  BCOUT(13) => R1IN_2_1_BCOUT(13),
  BCOUT(14) => R1IN_2_1_BCOUT(14),
  BCOUT(15) => R1IN_2_1_BCOUT(15),
  BCOUT(16) => R1IN_2_1_BCOUT(16),
  BCOUT(17) => R1IN_2_1_BCOUT(17),
  P(0) => R1IN_2F_0(0),
  P(1) => R1IN_2F_0(1),
  P(2) => R1IN_2F_0(2),
  P(3) => R1IN_2F_0(3),
  P(4) => R1IN_2F_0(4),
  P(5) => R1IN_2F_0(5),
  P(6) => R1IN_2F_0(6),
  P(7) => R1IN_2F_0(7),
  P(8) => R1IN_2F_0(8),
  P(9) => R1IN_2F_0(9),
  P(10) => R1IN_2F_0(10),
  P(11) => R1IN_2F_0(11),
  P(12) => R1IN_2F_0(12),
  P(13) => R1IN_2F_0(13),
  P(14) => R1IN_2F_0(14),
  P(15) => R1IN_2F_0(15),
  P(16) => R1IN_2F_0(16),
  P(17) => R1IN_2_1F_0(17),
  P(18) => R1IN_2_1F_0(18),
  P(19) => R1IN_2_1F_0(19),
  P(20) => R1IN_2_1F_0(20),
  P(21) => R1IN_2_1F_0(21),
  P(22) => R1IN_2_1F_0(22),
  P(23) => R1IN_2_1F_0(23),
  P(24) => R1IN_2_1F_0(24),
  P(25) => R1IN_2_1F_0(25),
  P(26) => R1IN_2_1F_0(26),
  P(27) => R1IN_2_1F_0(27),
  P(28) => R1IN_2_1F_0(28),
  P(29) => R1IN_2_1F_0(29),
  P(30) => R1IN_2_1F_0(30),
  P(31) => R1IN_2_1F_0(31),
  P(32) => R1IN_2_1F_0(32),
  P(33) => R1IN_2_1F_0(33),
  P(34) => UC_173_0,
  P(35) => UC_174_0,
  P(36) => UC_175_0,
  P(37) => UC_176_0,
  P(38) => UC_177_0,
  P(39) => UC_178_0,
  P(40) => UC_179_0,
  P(41) => UC_180_0,
  P(42) => UC_181_0,
  P(43) => UC_182_0,
  P(44) => UC_183_0,
  P(45) => UC_184_0,
  P(46) => UC_185_0,
  P(47) => UC_186_0,
  PCOUT(0) => R1IN_2_1_PCOUT(0),
  PCOUT(1) => R1IN_2_1_PCOUT(1),
  PCOUT(2) => R1IN_2_1_PCOUT(2),
  PCOUT(3) => R1IN_2_1_PCOUT(3),
  PCOUT(4) => R1IN_2_1_PCOUT(4),
  PCOUT(5) => R1IN_2_1_PCOUT(5),
  PCOUT(6) => R1IN_2_1_PCOUT(6),
  PCOUT(7) => R1IN_2_1_PCOUT(7),
  PCOUT(8) => R1IN_2_1_PCOUT(8),
  PCOUT(9) => R1IN_2_1_PCOUT(9),
  PCOUT(10) => R1IN_2_1_PCOUT(10),
  PCOUT(11) => R1IN_2_1_PCOUT(11),
  PCOUT(12) => R1IN_2_1_PCOUT(12),
  PCOUT(13) => R1IN_2_1_PCOUT(13),
  PCOUT(14) => R1IN_2_1_PCOUT(14),
  PCOUT(15) => R1IN_2_1_PCOUT(15),
  PCOUT(16) => R1IN_2_1_PCOUT(16),
  PCOUT(17) => R1IN_2_1_PCOUT(17),
  PCOUT(18) => R1IN_2_1_PCOUT(18),
  PCOUT(19) => R1IN_2_1_PCOUT(19),
  PCOUT(20) => R1IN_2_1_PCOUT(20),
  PCOUT(21) => R1IN_2_1_PCOUT(21),
  PCOUT(22) => R1IN_2_1_PCOUT(22),
  PCOUT(23) => R1IN_2_1_PCOUT(23),
  PCOUT(24) => R1IN_2_1_PCOUT(24),
  PCOUT(25) => R1IN_2_1_PCOUT(25),
  PCOUT(26) => R1IN_2_1_PCOUT(26),
  PCOUT(27) => R1IN_2_1_PCOUT(27),
  PCOUT(28) => R1IN_2_1_PCOUT(28),
  PCOUT(29) => R1IN_2_1_PCOUT(29),
  PCOUT(30) => R1IN_2_1_PCOUT(30),
  PCOUT(31) => R1IN_2_1_PCOUT(31),
  PCOUT(32) => R1IN_2_1_PCOUT(32),
  PCOUT(33) => R1IN_2_1_PCOUT(33),
  PCOUT(34) => R1IN_2_1_PCOUT(34),
  PCOUT(35) => R1IN_2_1_PCOUT(35),
  PCOUT(36) => R1IN_2_1_PCOUT(36),
  PCOUT(37) => R1IN_2_1_PCOUT(37),
  PCOUT(38) => R1IN_2_1_PCOUT(38),
  PCOUT(39) => R1IN_2_1_PCOUT(39),
  PCOUT(40) => R1IN_2_1_PCOUT(40),
  PCOUT(41) => R1IN_2_1_PCOUT(41),
  PCOUT(42) => R1IN_2_1_PCOUT(42),
  PCOUT(43) => R1IN_2_1_PCOUT(43),
  PCOUT(44) => R1IN_2_1_PCOUT(44),
  PCOUT(45) => R1IN_2_1_PCOUT(45),
  PCOUT(46) => R1IN_2_1_PCOUT(46),
  PCOUT(47) => R1IN_2_1_PCOUT(47));
\R1IN_1[33:0]\: DSP48 
generic map(
  AREG => 1,
  BREG => 1,
  CREG => 0,
  PREG => 1,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "CASCADE",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => A(0),
  A(1) => A(1),
  A(2) => A(2),
  A(3) => A(3),
  A(4) => A(4),
  A(5) => A(5),
  A(6) => A(6),
  A(7) => A(7),
  A(8) => A(8),
  A(9) => A(9),
  A(10) => A(10),
  A(11) => A(11),
  A(12) => A(12),
  A(13) => A(13),
  A(14) => A(14),
  A(15) => A(15),
  A(16) => A(16),
  A(17) => NN_1,
  B(0) => NN_1,
  B(1) => NN_1,
  B(2) => NN_1,
  B(3) => NN_1,
  B(4) => NN_1,
  B(5) => NN_1,
  B(6) => NN_1,
  B(7) => NN_1,
  B(8) => NN_1,
  B(9) => NN_1,
  B(10) => NN_1,
  B(11) => NN_1,
  B(12) => NN_1,
  B(13) => NN_1,
  B(14) => NN_1,
  B(15) => NN_1,
  B(16) => NN_1,
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => B_0(0),
  BCIN(1) => B_0(1),
  BCIN(2) => B_0(2),
  BCIN(3) => B_0(3),
  BCIN(4) => B_0(4),
  BCIN(5) => B_0(5),
  BCIN(6) => B_0(6),
  BCIN(7) => B_0(7),
  BCIN(8) => B_0(8),
  BCIN(9) => B_0(9),
  BCIN(10) => B_0(10),
  BCIN(11) => B_0(11),
  BCIN(12) => B_0(12),
  BCIN(13) => B_0(13),
  BCIN(14) => B_0(14),
  BCIN(15) => B_0(15),
  BCIN(16) => B_0(16),
  BCIN(17) => GND_0,
  PCIN(0) => NN_1,
  PCIN(1) => NN_1,
  PCIN(2) => NN_1,
  PCIN(3) => NN_1,
  PCIN(4) => NN_1,
  PCIN(5) => NN_1,
  PCIN(6) => NN_1,
  PCIN(7) => NN_1,
  PCIN(8) => NN_1,
  PCIN(9) => NN_1,
  PCIN(10) => NN_1,
  PCIN(11) => NN_1,
  PCIN(12) => NN_1,
  PCIN(13) => NN_1,
  PCIN(14) => NN_1,
  PCIN(15) => NN_1,
  PCIN(16) => NN_1,
  PCIN(17) => NN_1,
  PCIN(18) => NN_1,
  PCIN(19) => NN_1,
  PCIN(20) => NN_1,
  PCIN(21) => NN_1,
  PCIN(22) => NN_1,
  PCIN(23) => NN_1,
  PCIN(24) => NN_1,
  PCIN(25) => NN_1,
  PCIN(26) => NN_1,
  PCIN(27) => NN_1,
  PCIN(28) => NN_1,
  PCIN(29) => NN_1,
  PCIN(30) => NN_1,
  PCIN(31) => NN_1,
  PCIN(32) => NN_1,
  PCIN(33) => NN_1,
  PCIN(34) => NN_1,
  PCIN(35) => NN_1,
  PCIN(36) => NN_1,
  PCIN(37) => NN_1,
  PCIN(38) => NN_1,
  PCIN(39) => NN_1,
  PCIN(40) => NN_1,
  PCIN(41) => NN_1,
  PCIN(42) => NN_1,
  PCIN(43) => NN_1,
  PCIN(44) => NN_1,
  PCIN(45) => NN_1,
  PCIN(46) => NN_1,
  PCIN(47) => NN_1,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_1,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => CLK,
  CEA => EN,
  CEB => EN,
  CEC => NN_1,
  CEP => EN,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_1_BCOUT(0),
  BCOUT(1) => R1IN_1_BCOUT(1),
  BCOUT(2) => R1IN_1_BCOUT(2),
  BCOUT(3) => R1IN_1_BCOUT(3),
  BCOUT(4) => R1IN_1_BCOUT(4),
  BCOUT(5) => R1IN_1_BCOUT(5),
  BCOUT(6) => R1IN_1_BCOUT(6),
  BCOUT(7) => R1IN_1_BCOUT(7),
  BCOUT(8) => R1IN_1_BCOUT(8),
  BCOUT(9) => R1IN_1_BCOUT(9),
  BCOUT(10) => R1IN_1_BCOUT(10),
  BCOUT(11) => R1IN_1_BCOUT(11),
  BCOUT(12) => R1IN_1_BCOUT(12),
  BCOUT(13) => R1IN_1_BCOUT(13),
  BCOUT(14) => R1IN_1_BCOUT(14),
  BCOUT(15) => R1IN_1_BCOUT(15),
  BCOUT(16) => R1IN_1_BCOUT(16),
  BCOUT(17) => R1IN_1_BCOUT(17),
  P(0) => PRODUCT(0),
  P(1) => PRODUCT(1),
  P(2) => PRODUCT(2),
  P(3) => PRODUCT(3),
  P(4) => PRODUCT(4),
  P(5) => PRODUCT(5),
  P(6) => PRODUCT(6),
  P(7) => PRODUCT(7),
  P(8) => PRODUCT(8),
  P(9) => PRODUCT(9),
  P(10) => PRODUCT(10),
  P(11) => PRODUCT(11),
  P(12) => PRODUCT(12),
  P(13) => PRODUCT(13),
  P(14) => PRODUCT(14),
  P(15) => PRODUCT(15),
  P(16) => PRODUCT(16),
  P(17) => R1IN_ADD_2_0,
  P(18) => R1IN_1FF(18),
  P(19) => R1IN_1FF(19),
  P(20) => R1IN_1FF(20),
  P(21) => R1IN_1FF(21),
  P(22) => R1IN_1FF(22),
  P(23) => R1IN_1FF(23),
  P(24) => R1IN_1FF(24),
  P(25) => R1IN_1FF(25),
  P(26) => R1IN_1FF(26),
  P(27) => R1IN_1FF(27),
  P(28) => R1IN_1FF(28),
  P(29) => R1IN_1FF(29),
  P(30) => R1IN_1FF(30),
  P(31) => R1IN_1FF(31),
  P(32) => R1IN_1FF(32),
  P(33) => R1IN_1FF(33),
  P(34) => UC_159,
  P(35) => UC_160,
  P(36) => UC_161,
  P(37) => UC_162,
  P(38) => UC_163,
  P(39) => UC_164,
  P(40) => UC_165,
  P(41) => UC_166,
  P(42) => UC_167,
  P(43) => UC_168,
  P(44) => UC_169,
  P(45) => UC_170,
  P(46) => UC_171,
  P(47) => UC_172,
  PCOUT(0) => R1IN_1_PCOUT(0),
  PCOUT(1) => R1IN_1_PCOUT(1),
  PCOUT(2) => R1IN_1_PCOUT(2),
  PCOUT(3) => R1IN_1_PCOUT(3),
  PCOUT(4) => R1IN_1_PCOUT(4),
  PCOUT(5) => R1IN_1_PCOUT(5),
  PCOUT(6) => R1IN_1_PCOUT(6),
  PCOUT(7) => R1IN_1_PCOUT(7),
  PCOUT(8) => R1IN_1_PCOUT(8),
  PCOUT(9) => R1IN_1_PCOUT(9),
  PCOUT(10) => R1IN_1_PCOUT(10),
  PCOUT(11) => R1IN_1_PCOUT(11),
  PCOUT(12) => R1IN_1_PCOUT(12),
  PCOUT(13) => R1IN_1_PCOUT(13),
  PCOUT(14) => R1IN_1_PCOUT(14),
  PCOUT(15) => R1IN_1_PCOUT(15),
  PCOUT(16) => R1IN_1_PCOUT(16),
  PCOUT(17) => R1IN_1_PCOUT(17),
  PCOUT(18) => R1IN_1_PCOUT(18),
  PCOUT(19) => R1IN_1_PCOUT(19),
  PCOUT(20) => R1IN_1_PCOUT(20),
  PCOUT(21) => R1IN_1_PCOUT(21),
  PCOUT(22) => R1IN_1_PCOUT(22),
  PCOUT(23) => R1IN_1_PCOUT(23),
  PCOUT(24) => R1IN_1_PCOUT(24),
  PCOUT(25) => R1IN_1_PCOUT(25),
  PCOUT(26) => R1IN_1_PCOUT(26),
  PCOUT(27) => R1IN_1_PCOUT(27),
  PCOUT(28) => R1IN_1_PCOUT(28),
  PCOUT(29) => R1IN_1_PCOUT(29),
  PCOUT(30) => R1IN_1_PCOUT(30),
  PCOUT(31) => R1IN_1_PCOUT(31),
  PCOUT(32) => R1IN_1_PCOUT(32),
  PCOUT(33) => R1IN_1_PCOUT(33),
  PCOUT(34) => R1IN_1_PCOUT(34),
  PCOUT(35) => R1IN_1_PCOUT(35),
  PCOUT(36) => R1IN_1_PCOUT(36),
  PCOUT(37) => R1IN_1_PCOUT(37),
  PCOUT(38) => R1IN_1_PCOUT(38),
  PCOUT(39) => R1IN_1_PCOUT(39),
  PCOUT(40) => R1IN_1_PCOUT(40),
  PCOUT(41) => R1IN_1_PCOUT(41),
  PCOUT(42) => R1IN_1_PCOUT(42),
  PCOUT(43) => R1IN_1_PCOUT(43),
  PCOUT(44) => R1IN_1_PCOUT(44),
  PCOUT(45) => R1IN_1_PCOUT(45),
  PCOUT(46) => R1IN_1_PCOUT(46),
  PCOUT(47) => R1IN_1_PCOUT(47));
\R1IN_4_3_1[33:0]\: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 0,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => B(34),
  A(1) => B(35),
  A(2) => B(36),
  A(3) => B(37),
  A(4) => B(38),
  A(5) => B(39),
  A(6) => B(40),
  A(7) => B(41),
  A(8) => B(42),
  A(9) => B(43),
  A(10) => B(44),
  A(11) => B(45),
  A(12) => B(46),
  A(13) => B(47),
  A(14) => B(48),
  A(15) => B(49),
  A(16) => B(50),
  A(17) => NN_1,
  B(0) => A(17),
  B(1) => A(18),
  B(2) => A(19),
  B(3) => A(20),
  B(4) => A(21),
  B(5) => A(22),
  B(6) => A(23),
  B(7) => A(24),
  B(8) => A(25),
  B(9) => A(26),
  B(10) => A(27),
  B(11) => A(28),
  B(12) => A(29),
  B(13) => A(30),
  B(14) => A(31),
  B(15) => A(32),
  B(16) => A(33),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => NN_1,
  PCIN(1) => NN_1,
  PCIN(2) => NN_1,
  PCIN(3) => NN_1,
  PCIN(4) => NN_1,
  PCIN(5) => NN_1,
  PCIN(6) => NN_1,
  PCIN(7) => NN_1,
  PCIN(8) => NN_1,
  PCIN(9) => NN_1,
  PCIN(10) => NN_1,
  PCIN(11) => NN_1,
  PCIN(12) => NN_1,
  PCIN(13) => NN_1,
  PCIN(14) => NN_1,
  PCIN(15) => NN_1,
  PCIN(16) => NN_1,
  PCIN(17) => NN_1,
  PCIN(18) => NN_1,
  PCIN(19) => NN_1,
  PCIN(20) => NN_1,
  PCIN(21) => NN_1,
  PCIN(22) => NN_1,
  PCIN(23) => NN_1,
  PCIN(24) => NN_1,
  PCIN(25) => NN_1,
  PCIN(26) => NN_1,
  PCIN(27) => NN_1,
  PCIN(28) => NN_1,
  PCIN(29) => NN_1,
  PCIN(30) => NN_1,
  PCIN(31) => NN_1,
  PCIN(32) => NN_1,
  PCIN(33) => NN_1,
  PCIN(34) => NN_1,
  PCIN(35) => NN_1,
  PCIN(36) => NN_1,
  PCIN(37) => NN_1,
  PCIN(38) => NN_1,
  PCIN(39) => NN_1,
  PCIN(40) => NN_1,
  PCIN(41) => NN_1,
  PCIN(42) => NN_1,
  PCIN(43) => NN_1,
  PCIN(44) => NN_1,
  PCIN(45) => NN_1,
  PCIN(46) => NN_1,
  PCIN(47) => NN_1,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_1,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => NN_1,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => NN_1,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_4_3_1_BCOUT(0),
  BCOUT(1) => R1IN_4_3_1_BCOUT(1),
  BCOUT(2) => R1IN_4_3_1_BCOUT(2),
  BCOUT(3) => R1IN_4_3_1_BCOUT(3),
  BCOUT(4) => R1IN_4_3_1_BCOUT(4),
  BCOUT(5) => R1IN_4_3_1_BCOUT(5),
  BCOUT(6) => R1IN_4_3_1_BCOUT(6),
  BCOUT(7) => R1IN_4_3_1_BCOUT(7),
  BCOUT(8) => R1IN_4_3_1_BCOUT(8),
  BCOUT(9) => R1IN_4_3_1_BCOUT(9),
  BCOUT(10) => R1IN_4_3_1_BCOUT(10),
  BCOUT(11) => R1IN_4_3_1_BCOUT(11),
  BCOUT(12) => R1IN_4_3_1_BCOUT(12),
  BCOUT(13) => R1IN_4_3_1_BCOUT(13),
  BCOUT(14) => R1IN_4_3_1_BCOUT(14),
  BCOUT(15) => R1IN_4_3_1_BCOUT(15),
  BCOUT(16) => R1IN_4_3_1_BCOUT(16),
  BCOUT(17) => R1IN_4_3_1_BCOUT(17),
  P(0) => R1IN_4_3(0),
  P(1) => R1IN_4_3(1),
  P(2) => R1IN_4_3(2),
  P(3) => R1IN_4_3(3),
  P(4) => R1IN_4_3(4),
  P(5) => R1IN_4_3(5),
  P(6) => R1IN_4_3(6),
  P(7) => R1IN_4_3(7),
  P(8) => R1IN_4_3(8),
  P(9) => R1IN_4_3(9),
  P(10) => R1IN_4_3(10),
  P(11) => R1IN_4_3(11),
  P(12) => R1IN_4_3(12),
  P(13) => R1IN_4_3(13),
  P(14) => R1IN_4_3(14),
  P(15) => R1IN_4_3(15),
  P(16) => R1IN_4_3(16),
  P(17) => R1IN_4_3_1(17),
  P(18) => R1IN_4_3_1(18),
  P(19) => R1IN_4_3_1(19),
  P(20) => R1IN_4_3_1(20),
  P(21) => R1IN_4_3_1(21),
  P(22) => R1IN_4_3_1(22),
  P(23) => R1IN_4_3_1(23),
  P(24) => R1IN_4_3_1(24),
  P(25) => R1IN_4_3_1(25),
  P(26) => R1IN_4_3_1(26),
  P(27) => R1IN_4_3_1(27),
  P(28) => R1IN_4_3_1(28),
  P(29) => R1IN_4_3_1(29),
  P(30) => R1IN_4_3_1(30),
  P(31) => R1IN_4_3_1(31),
  P(32) => R1IN_4_3_1(32),
  P(33) => R1IN_4_3_1(33),
  P(34) => UC_145,
  P(35) => UC_146,
  P(36) => UC_147,
  P(37) => UC_148,
  P(38) => UC_149,
  P(39) => UC_150,
  P(40) => UC_151,
  P(41) => UC_152,
  P(42) => UC_153,
  P(43) => UC_154,
  P(44) => UC_155,
  P(45) => UC_156,
  P(46) => UC_157,
  P(47) => UC_158,
  PCOUT(0) => R1IN_4_3_0(0),
  PCOUT(1) => R1IN_4_3_0(1),
  PCOUT(2) => R1IN_4_3_0(2),
  PCOUT(3) => R1IN_4_3_0(3),
  PCOUT(4) => R1IN_4_3_0(4),
  PCOUT(5) => R1IN_4_3_0(5),
  PCOUT(6) => R1IN_4_3_0(6),
  PCOUT(7) => R1IN_4_3_0(7),
  PCOUT(8) => R1IN_4_3_0(8),
  PCOUT(9) => R1IN_4_3_0(9),
  PCOUT(10) => R1IN_4_3_0(10),
  PCOUT(11) => R1IN_4_3_0(11),
  PCOUT(12) => R1IN_4_3_0(12),
  PCOUT(13) => R1IN_4_3_0(13),
  PCOUT(14) => R1IN_4_3_0(14),
  PCOUT(15) => R1IN_4_3_0(15),
  PCOUT(16) => R1IN_4_3_0(16),
  PCOUT(17) => R1IN_4_3_1_0(17),
  PCOUT(18) => R1IN_4_3_1_0(18),
  PCOUT(19) => R1IN_4_3_1_0(19),
  PCOUT(20) => R1IN_4_3_1_0(20),
  PCOUT(21) => R1IN_4_3_1_0(21),
  PCOUT(22) => R1IN_4_3_1_0(22),
  PCOUT(23) => R1IN_4_3_1_0(23),
  PCOUT(24) => R1IN_4_3_1_0(24),
  PCOUT(25) => R1IN_4_3_1_0(25),
  PCOUT(26) => R1IN_4_3_1_0(26),
  PCOUT(27) => R1IN_4_3_1_0(27),
  PCOUT(28) => R1IN_4_3_1_0(28),
  PCOUT(29) => R1IN_4_3_1_0(29),
  PCOUT(30) => R1IN_4_3_1_0(30),
  PCOUT(31) => R1IN_4_3_1_0(31),
  PCOUT(32) => R1IN_4_3_1_0(32),
  PCOUT(33) => R1IN_4_3_1_0(33),
  PCOUT(34) => UC_145_0,
  PCOUT(35) => UC_146_0,
  PCOUT(36) => UC_147_0,
  PCOUT(37) => UC_148_0,
  PCOUT(38) => UC_149_0,
  PCOUT(39) => UC_150_0,
  PCOUT(40) => UC_151_0,
  PCOUT(41) => UC_152_0,
  PCOUT(42) => UC_153_0,
  PCOUT(43) => UC_154_0,
  PCOUT(44) => UC_155_0,
  PCOUT(45) => UC_156_0,
  PCOUT(46) => UC_157_0,
  PCOUT(47) => UC_158_0);
\R1IN_4_2_1[33:0]\: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 0,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => A(34),
  A(1) => A(35),
  A(2) => A(36),
  A(3) => A(37),
  A(4) => A(38),
  A(5) => A(39),
  A(6) => A(40),
  A(7) => A(41),
  A(8) => A(42),
  A(9) => A(43),
  A(10) => A(44),
  A(11) => A(45),
  A(12) => A(46),
  A(13) => A(47),
  A(14) => A(48),
  A(15) => A(49),
  A(16) => A(50),
  A(17) => NN_1,
  B(0) => B(17),
  B(1) => B(18),
  B(2) => B(19),
  B(3) => B(20),
  B(4) => B(21),
  B(5) => B(22),
  B(6) => B(23),
  B(7) => B(24),
  B(8) => B(25),
  B(9) => B(26),
  B(10) => B(27),
  B(11) => B(28),
  B(12) => B(29),
  B(13) => B(30),
  B(14) => B(31),
  B(15) => B(32),
  B(16) => B(33),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => NN_1,
  PCIN(1) => NN_1,
  PCIN(2) => NN_1,
  PCIN(3) => NN_1,
  PCIN(4) => NN_1,
  PCIN(5) => NN_1,
  PCIN(6) => NN_1,
  PCIN(7) => NN_1,
  PCIN(8) => NN_1,
  PCIN(9) => NN_1,
  PCIN(10) => NN_1,
  PCIN(11) => NN_1,
  PCIN(12) => NN_1,
  PCIN(13) => NN_1,
  PCIN(14) => NN_1,
  PCIN(15) => NN_1,
  PCIN(16) => NN_1,
  PCIN(17) => NN_1,
  PCIN(18) => NN_1,
  PCIN(19) => NN_1,
  PCIN(20) => NN_1,
  PCIN(21) => NN_1,
  PCIN(22) => NN_1,
  PCIN(23) => NN_1,
  PCIN(24) => NN_1,
  PCIN(25) => NN_1,
  PCIN(26) => NN_1,
  PCIN(27) => NN_1,
  PCIN(28) => NN_1,
  PCIN(29) => NN_1,
  PCIN(30) => NN_1,
  PCIN(31) => NN_1,
  PCIN(32) => NN_1,
  PCIN(33) => NN_1,
  PCIN(34) => NN_1,
  PCIN(35) => NN_1,
  PCIN(36) => NN_1,
  PCIN(37) => NN_1,
  PCIN(38) => NN_1,
  PCIN(39) => NN_1,
  PCIN(40) => NN_1,
  PCIN(41) => NN_1,
  PCIN(42) => NN_1,
  PCIN(43) => NN_1,
  PCIN(44) => NN_1,
  PCIN(45) => NN_1,
  PCIN(46) => NN_1,
  PCIN(47) => NN_1,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_1,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => NN_1,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => NN_1,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_4_2_1_BCOUT(0),
  BCOUT(1) => R1IN_4_2_1_BCOUT(1),
  BCOUT(2) => R1IN_4_2_1_BCOUT(2),
  BCOUT(3) => R1IN_4_2_1_BCOUT(3),
  BCOUT(4) => R1IN_4_2_1_BCOUT(4),
  BCOUT(5) => R1IN_4_2_1_BCOUT(5),
  BCOUT(6) => R1IN_4_2_1_BCOUT(6),
  BCOUT(7) => R1IN_4_2_1_BCOUT(7),
  BCOUT(8) => R1IN_4_2_1_BCOUT(8),
  BCOUT(9) => R1IN_4_2_1_BCOUT(9),
  BCOUT(10) => R1IN_4_2_1_BCOUT(10),
  BCOUT(11) => R1IN_4_2_1_BCOUT(11),
  BCOUT(12) => R1IN_4_2_1_BCOUT(12),
  BCOUT(13) => R1IN_4_2_1_BCOUT(13),
  BCOUT(14) => R1IN_4_2_1_BCOUT(14),
  BCOUT(15) => R1IN_4_2_1_BCOUT(15),
  BCOUT(16) => R1IN_4_2_1_BCOUT(16),
  BCOUT(17) => R1IN_4_2_1_BCOUT(17),
  P(0) => R1IN_4_2(0),
  P(1) => R1IN_4_2(1),
  P(2) => R1IN_4_2(2),
  P(3) => R1IN_4_2(3),
  P(4) => R1IN_4_2(4),
  P(5) => R1IN_4_2(5),
  P(6) => R1IN_4_2(6),
  P(7) => R1IN_4_2(7),
  P(8) => R1IN_4_2(8),
  P(9) => R1IN_4_2(9),
  P(10) => R1IN_4_2(10),
  P(11) => R1IN_4_2(11),
  P(12) => R1IN_4_2(12),
  P(13) => R1IN_4_2(13),
  P(14) => R1IN_4_2(14),
  P(15) => R1IN_4_2(15),
  P(16) => R1IN_4_2(16),
  P(17) => R1IN_4_2_1(17),
  P(18) => R1IN_4_2_1(18),
  P(19) => R1IN_4_2_1(19),
  P(20) => R1IN_4_2_1(20),
  P(21) => R1IN_4_2_1(21),
  P(22) => R1IN_4_2_1(22),
  P(23) => R1IN_4_2_1(23),
  P(24) => R1IN_4_2_1(24),
  P(25) => R1IN_4_2_1(25),
  P(26) => R1IN_4_2_1(26),
  P(27) => R1IN_4_2_1(27),
  P(28) => R1IN_4_2_1(28),
  P(29) => R1IN_4_2_1(29),
  P(30) => R1IN_4_2_1(30),
  P(31) => R1IN_4_2_1(31),
  P(32) => R1IN_4_2_1(32),
  P(33) => R1IN_4_2_1(33),
  P(34) => UC_131,
  P(35) => UC_132,
  P(36) => UC_133,
  P(37) => UC_134,
  P(38) => UC_135,
  P(39) => UC_136,
  P(40) => UC_137,
  P(41) => UC_138,
  P(42) => UC_139,
  P(43) => UC_140,
  P(44) => UC_141,
  P(45) => UC_142,
  P(46) => UC_143,
  P(47) => UC_144,
  PCOUT(0) => R1IN_4_2_0(0),
  PCOUT(1) => R1IN_4_2_0(1),
  PCOUT(2) => R1IN_4_2_0(2),
  PCOUT(3) => R1IN_4_2_0(3),
  PCOUT(4) => R1IN_4_2_0(4),
  PCOUT(5) => R1IN_4_2_0(5),
  PCOUT(6) => R1IN_4_2_0(6),
  PCOUT(7) => R1IN_4_2_0(7),
  PCOUT(8) => R1IN_4_2_0(8),
  PCOUT(9) => R1IN_4_2_0(9),
  PCOUT(10) => R1IN_4_2_0(10),
  PCOUT(11) => R1IN_4_2_0(11),
  PCOUT(12) => R1IN_4_2_0(12),
  PCOUT(13) => R1IN_4_2_0(13),
  PCOUT(14) => R1IN_4_2_0(14),
  PCOUT(15) => R1IN_4_2_0(15),
  PCOUT(16) => R1IN_4_2_0(16),
  PCOUT(17) => R1IN_4_2_1_0(17),
  PCOUT(18) => R1IN_4_2_1_0(18),
  PCOUT(19) => R1IN_4_2_1_0(19),
  PCOUT(20) => R1IN_4_2_1_0(20),
  PCOUT(21) => R1IN_4_2_1_0(21),
  PCOUT(22) => R1IN_4_2_1_0(22),
  PCOUT(23) => R1IN_4_2_1_0(23),
  PCOUT(24) => R1IN_4_2_1_0(24),
  PCOUT(25) => R1IN_4_2_1_0(25),
  PCOUT(26) => R1IN_4_2_1_0(26),
  PCOUT(27) => R1IN_4_2_1_0(27),
  PCOUT(28) => R1IN_4_2_1_0(28),
  PCOUT(29) => R1IN_4_2_1_0(29),
  PCOUT(30) => R1IN_4_2_1_0(30),
  PCOUT(31) => R1IN_4_2_1_0(31),
  PCOUT(32) => R1IN_4_2_1_0(32),
  PCOUT(33) => R1IN_4_2_1_0(33),
  PCOUT(34) => UC_131_0,
  PCOUT(35) => UC_132_0,
  PCOUT(36) => UC_133_0,
  PCOUT(37) => UC_134_0,
  PCOUT(38) => UC_135_0,
  PCOUT(39) => UC_136_0,
  PCOUT(40) => UC_137_0,
  PCOUT(41) => UC_138_0,
  PCOUT(42) => UC_139_0,
  PCOUT(43) => UC_140_0,
  PCOUT(44) => UC_141_0,
  PCOUT(45) => UC_142_0,
  PCOUT(46) => UC_143_0,
  PCOUT(47) => UC_144_0);
\R1IN_3_2_1[33:0]\: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 0,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => B(34),
  A(1) => B(35),
  A(2) => B(36),
  A(3) => B(37),
  A(4) => B(38),
  A(5) => B(39),
  A(6) => B(40),
  A(7) => B(41),
  A(8) => B(42),
  A(9) => B(43),
  A(10) => B(44),
  A(11) => B(45),
  A(12) => B(46),
  A(13) => B(47),
  A(14) => B(48),
  A(15) => B(49),
  A(16) => B(50),
  A(17) => NN_1,
  B(0) => A(0),
  B(1) => A(1),
  B(2) => A(2),
  B(3) => A(3),
  B(4) => A(4),
  B(5) => A(5),
  B(6) => A(6),
  B(7) => A(7),
  B(8) => A(8),
  B(9) => A(9),
  B(10) => A(10),
  B(11) => A(11),
  B(12) => A(12),
  B(13) => A(13),
  B(14) => A(14),
  B(15) => A(15),
  B(16) => A(16),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => NN_1,
  PCIN(1) => NN_1,
  PCIN(2) => NN_1,
  PCIN(3) => NN_1,
  PCIN(4) => NN_1,
  PCIN(5) => NN_1,
  PCIN(6) => NN_1,
  PCIN(7) => NN_1,
  PCIN(8) => NN_1,
  PCIN(9) => NN_1,
  PCIN(10) => NN_1,
  PCIN(11) => NN_1,
  PCIN(12) => NN_1,
  PCIN(13) => NN_1,
  PCIN(14) => NN_1,
  PCIN(15) => NN_1,
  PCIN(16) => NN_1,
  PCIN(17) => NN_1,
  PCIN(18) => NN_1,
  PCIN(19) => NN_1,
  PCIN(20) => NN_1,
  PCIN(21) => NN_1,
  PCIN(22) => NN_1,
  PCIN(23) => NN_1,
  PCIN(24) => NN_1,
  PCIN(25) => NN_1,
  PCIN(26) => NN_1,
  PCIN(27) => NN_1,
  PCIN(28) => NN_1,
  PCIN(29) => NN_1,
  PCIN(30) => NN_1,
  PCIN(31) => NN_1,
  PCIN(32) => NN_1,
  PCIN(33) => NN_1,
  PCIN(34) => NN_1,
  PCIN(35) => NN_1,
  PCIN(36) => NN_1,
  PCIN(37) => NN_1,
  PCIN(38) => NN_1,
  PCIN(39) => NN_1,
  PCIN(40) => NN_1,
  PCIN(41) => NN_1,
  PCIN(42) => NN_1,
  PCIN(43) => NN_1,
  PCIN(44) => NN_1,
  PCIN(45) => NN_1,
  PCIN(46) => NN_1,
  PCIN(47) => NN_1,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_1,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => NN_1,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => NN_1,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_3_2_1_BCOUT(0),
  BCOUT(1) => R1IN_3_2_1_BCOUT(1),
  BCOUT(2) => R1IN_3_2_1_BCOUT(2),
  BCOUT(3) => R1IN_3_2_1_BCOUT(3),
  BCOUT(4) => R1IN_3_2_1_BCOUT(4),
  BCOUT(5) => R1IN_3_2_1_BCOUT(5),
  BCOUT(6) => R1IN_3_2_1_BCOUT(6),
  BCOUT(7) => R1IN_3_2_1_BCOUT(7),
  BCOUT(8) => R1IN_3_2_1_BCOUT(8),
  BCOUT(9) => R1IN_3_2_1_BCOUT(9),
  BCOUT(10) => R1IN_3_2_1_BCOUT(10),
  BCOUT(11) => R1IN_3_2_1_BCOUT(11),
  BCOUT(12) => R1IN_3_2_1_BCOUT(12),
  BCOUT(13) => R1IN_3_2_1_BCOUT(13),
  BCOUT(14) => R1IN_3_2_1_BCOUT(14),
  BCOUT(15) => R1IN_3_2_1_BCOUT(15),
  BCOUT(16) => R1IN_3_2_1_BCOUT(16),
  BCOUT(17) => R1IN_3_2_1_BCOUT(17),
  P(0) => R1IN_3_2(0),
  P(1) => R1IN_3_2(1),
  P(2) => R1IN_3_2(2),
  P(3) => R1IN_3_2(3),
  P(4) => R1IN_3_2(4),
  P(5) => R1IN_3_2(5),
  P(6) => R1IN_3_2(6),
  P(7) => R1IN_3_2(7),
  P(8) => R1IN_3_2(8),
  P(9) => R1IN_3_2(9),
  P(10) => R1IN_3_2(10),
  P(11) => R1IN_3_2(11),
  P(12) => R1IN_3_2(12),
  P(13) => R1IN_3_2(13),
  P(14) => R1IN_3_2(14),
  P(15) => R1IN_3_2(15),
  P(16) => R1IN_3_2(16),
  P(17) => R1IN_3_2_1(17),
  P(18) => R1IN_3_2_1(18),
  P(19) => R1IN_3_2_1(19),
  P(20) => R1IN_3_2_1(20),
  P(21) => R1IN_3_2_1(21),
  P(22) => R1IN_3_2_1(22),
  P(23) => R1IN_3_2_1(23),
  P(24) => R1IN_3_2_1(24),
  P(25) => R1IN_3_2_1(25),
  P(26) => R1IN_3_2_1(26),
  P(27) => R1IN_3_2_1(27),
  P(28) => R1IN_3_2_1(28),
  P(29) => R1IN_3_2_1(29),
  P(30) => R1IN_3_2_1(30),
  P(31) => R1IN_3_2_1(31),
  P(32) => R1IN_3_2_1(32),
  P(33) => R1IN_3_2_1(33),
  P(34) => UC_117,
  P(35) => UC_118,
  P(36) => UC_119,
  P(37) => UC_120,
  P(38) => UC_121,
  P(39) => UC_122,
  P(40) => UC_123,
  P(41) => UC_124,
  P(42) => UC_125,
  P(43) => UC_126,
  P(44) => UC_127,
  P(45) => UC_128,
  P(46) => UC_129,
  P(47) => UC_130,
  PCOUT(0) => R1IN_3_2_0(0),
  PCOUT(1) => R1IN_3_2_0(1),
  PCOUT(2) => R1IN_3_2_0(2),
  PCOUT(3) => R1IN_3_2_0(3),
  PCOUT(4) => R1IN_3_2_0(4),
  PCOUT(5) => R1IN_3_2_0(5),
  PCOUT(6) => R1IN_3_2_0(6),
  PCOUT(7) => R1IN_3_2_0(7),
  PCOUT(8) => R1IN_3_2_0(8),
  PCOUT(9) => R1IN_3_2_0(9),
  PCOUT(10) => R1IN_3_2_0(10),
  PCOUT(11) => R1IN_3_2_0(11),
  PCOUT(12) => R1IN_3_2_0(12),
  PCOUT(13) => R1IN_3_2_0(13),
  PCOUT(14) => R1IN_3_2_0(14),
  PCOUT(15) => R1IN_3_2_0(15),
  PCOUT(16) => R1IN_3_2_0(16),
  PCOUT(17) => R1IN_3_2_1_0(17),
  PCOUT(18) => R1IN_3_2_1_0(18),
  PCOUT(19) => R1IN_3_2_1_0(19),
  PCOUT(20) => R1IN_3_2_1_0(20),
  PCOUT(21) => R1IN_3_2_1_0(21),
  PCOUT(22) => R1IN_3_2_1_0(22),
  PCOUT(23) => R1IN_3_2_1_0(23),
  PCOUT(24) => R1IN_3_2_1_0(24),
  PCOUT(25) => R1IN_3_2_1_0(25),
  PCOUT(26) => R1IN_3_2_1_0(26),
  PCOUT(27) => R1IN_3_2_1_0(27),
  PCOUT(28) => R1IN_3_2_1_0(28),
  PCOUT(29) => R1IN_3_2_1_0(29),
  PCOUT(30) => R1IN_3_2_1_0(30),
  PCOUT(31) => R1IN_3_2_1_0(31),
  PCOUT(32) => R1IN_3_2_1_0(32),
  PCOUT(33) => R1IN_3_2_1_0(33),
  PCOUT(34) => UC_117_0,
  PCOUT(35) => UC_118_0,
  PCOUT(36) => UC_119_0,
  PCOUT(37) => UC_120_0,
  PCOUT(38) => UC_121_0,
  PCOUT(39) => UC_122_0,
  PCOUT(40) => UC_123_0,
  PCOUT(41) => UC_124_0,
  PCOUT(42) => UC_125_0,
  PCOUT(43) => UC_126_0,
  PCOUT(44) => UC_127_0,
  PCOUT(45) => UC_128_0,
  PCOUT(46) => UC_129_0,
  PCOUT(47) => UC_130_0);
\R1IN_2_2_1[33:0]\: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 0,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => A(34),
  A(1) => A(35),
  A(2) => A(36),
  A(3) => A(37),
  A(4) => A(38),
  A(5) => A(39),
  A(6) => A(40),
  A(7) => A(41),
  A(8) => A(42),
  A(9) => A(43),
  A(10) => A(44),
  A(11) => A(45),
  A(12) => A(46),
  A(13) => A(47),
  A(14) => A(48),
  A(15) => A(49),
  A(16) => A(50),
  A(17) => NN_1,
  B(0) => B(0),
  B(1) => B(1),
  B(2) => B(2),
  B(3) => B(3),
  B(4) => B(4),
  B(5) => B(5),
  B(6) => B(6),
  B(7) => B(7),
  B(8) => B(8),
  B(9) => B(9),
  B(10) => B(10),
  B(11) => B(11),
  B(12) => B(12),
  B(13) => B(13),
  B(14) => B(14),
  B(15) => B(15),
  B(16) => B(16),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => NN_1,
  PCIN(1) => NN_1,
  PCIN(2) => NN_1,
  PCIN(3) => NN_1,
  PCIN(4) => NN_1,
  PCIN(5) => NN_1,
  PCIN(6) => NN_1,
  PCIN(7) => NN_1,
  PCIN(8) => NN_1,
  PCIN(9) => NN_1,
  PCIN(10) => NN_1,
  PCIN(11) => NN_1,
  PCIN(12) => NN_1,
  PCIN(13) => NN_1,
  PCIN(14) => NN_1,
  PCIN(15) => NN_1,
  PCIN(16) => NN_1,
  PCIN(17) => NN_1,
  PCIN(18) => NN_1,
  PCIN(19) => NN_1,
  PCIN(20) => NN_1,
  PCIN(21) => NN_1,
  PCIN(22) => NN_1,
  PCIN(23) => NN_1,
  PCIN(24) => NN_1,
  PCIN(25) => NN_1,
  PCIN(26) => NN_1,
  PCIN(27) => NN_1,
  PCIN(28) => NN_1,
  PCIN(29) => NN_1,
  PCIN(30) => NN_1,
  PCIN(31) => NN_1,
  PCIN(32) => NN_1,
  PCIN(33) => NN_1,
  PCIN(34) => NN_1,
  PCIN(35) => NN_1,
  PCIN(36) => NN_1,
  PCIN(37) => NN_1,
  PCIN(38) => NN_1,
  PCIN(39) => NN_1,
  PCIN(40) => NN_1,
  PCIN(41) => NN_1,
  PCIN(42) => NN_1,
  PCIN(43) => NN_1,
  PCIN(44) => NN_1,
  PCIN(45) => NN_1,
  PCIN(46) => NN_1,
  PCIN(47) => NN_1,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_1,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => NN_1,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => NN_1,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_2_2_1_BCOUT(0),
  BCOUT(1) => R1IN_2_2_1_BCOUT(1),
  BCOUT(2) => R1IN_2_2_1_BCOUT(2),
  BCOUT(3) => R1IN_2_2_1_BCOUT(3),
  BCOUT(4) => R1IN_2_2_1_BCOUT(4),
  BCOUT(5) => R1IN_2_2_1_BCOUT(5),
  BCOUT(6) => R1IN_2_2_1_BCOUT(6),
  BCOUT(7) => R1IN_2_2_1_BCOUT(7),
  BCOUT(8) => R1IN_2_2_1_BCOUT(8),
  BCOUT(9) => R1IN_2_2_1_BCOUT(9),
  BCOUT(10) => R1IN_2_2_1_BCOUT(10),
  BCOUT(11) => R1IN_2_2_1_BCOUT(11),
  BCOUT(12) => R1IN_2_2_1_BCOUT(12),
  BCOUT(13) => R1IN_2_2_1_BCOUT(13),
  BCOUT(14) => R1IN_2_2_1_BCOUT(14),
  BCOUT(15) => R1IN_2_2_1_BCOUT(15),
  BCOUT(16) => R1IN_2_2_1_BCOUT(16),
  BCOUT(17) => R1IN_2_2_1_BCOUT(17),
  P(0) => R1IN_2_2(0),
  P(1) => R1IN_2_2(1),
  P(2) => R1IN_2_2(2),
  P(3) => R1IN_2_2(3),
  P(4) => R1IN_2_2(4),
  P(5) => R1IN_2_2(5),
  P(6) => R1IN_2_2(6),
  P(7) => R1IN_2_2(7),
  P(8) => R1IN_2_2(8),
  P(9) => R1IN_2_2(9),
  P(10) => R1IN_2_2(10),
  P(11) => R1IN_2_2(11),
  P(12) => R1IN_2_2(12),
  P(13) => R1IN_2_2(13),
  P(14) => R1IN_2_2(14),
  P(15) => R1IN_2_2(15),
  P(16) => R1IN_2_2(16),
  P(17) => R1IN_2_2_1(17),
  P(18) => R1IN_2_2_1(18),
  P(19) => R1IN_2_2_1(19),
  P(20) => R1IN_2_2_1(20),
  P(21) => R1IN_2_2_1(21),
  P(22) => R1IN_2_2_1(22),
  P(23) => R1IN_2_2_1(23),
  P(24) => R1IN_2_2_1(24),
  P(25) => R1IN_2_2_1(25),
  P(26) => R1IN_2_2_1(26),
  P(27) => R1IN_2_2_1(27),
  P(28) => R1IN_2_2_1(28),
  P(29) => R1IN_2_2_1(29),
  P(30) => R1IN_2_2_1(30),
  P(31) => R1IN_2_2_1(31),
  P(32) => R1IN_2_2_1(32),
  P(33) => R1IN_2_2_1(33),
  P(34) => UC_103,
  P(35) => UC_104,
  P(36) => UC_105,
  P(37) => UC_106,
  P(38) => UC_107,
  P(39) => UC_108,
  P(40) => UC_109,
  P(41) => UC_110,
  P(42) => UC_111,
  P(43) => UC_112,
  P(44) => UC_113,
  P(45) => UC_114,
  P(46) => UC_115,
  P(47) => UC_116,
  PCOUT(0) => R1IN_2_2_0(0),
  PCOUT(1) => R1IN_2_2_0(1),
  PCOUT(2) => R1IN_2_2_0(2),
  PCOUT(3) => R1IN_2_2_0(3),
  PCOUT(4) => R1IN_2_2_0(4),
  PCOUT(5) => R1IN_2_2_0(5),
  PCOUT(6) => R1IN_2_2_0(6),
  PCOUT(7) => R1IN_2_2_0(7),
  PCOUT(8) => R1IN_2_2_0(8),
  PCOUT(9) => R1IN_2_2_0(9),
  PCOUT(10) => R1IN_2_2_0(10),
  PCOUT(11) => R1IN_2_2_0(11),
  PCOUT(12) => R1IN_2_2_0(12),
  PCOUT(13) => R1IN_2_2_0(13),
  PCOUT(14) => R1IN_2_2_0(14),
  PCOUT(15) => R1IN_2_2_0(15),
  PCOUT(16) => R1IN_2_2_0(16),
  PCOUT(17) => R1IN_2_2_1_0(17),
  PCOUT(18) => R1IN_2_2_1_0(18),
  PCOUT(19) => R1IN_2_2_1_0(19),
  PCOUT(20) => R1IN_2_2_1_0(20),
  PCOUT(21) => R1IN_2_2_1_0(21),
  PCOUT(22) => R1IN_2_2_1_0(22),
  PCOUT(23) => R1IN_2_2_1_0(23),
  PCOUT(24) => R1IN_2_2_1_0(24),
  PCOUT(25) => R1IN_2_2_1_0(25),
  PCOUT(26) => R1IN_2_2_1_0(26),
  PCOUT(27) => R1IN_2_2_1_0(27),
  PCOUT(28) => R1IN_2_2_1_0(28),
  PCOUT(29) => R1IN_2_2_1_0(29),
  PCOUT(30) => R1IN_2_2_1_0(30),
  PCOUT(31) => R1IN_2_2_1_0(31),
  PCOUT(32) => R1IN_2_2_1_0(32),
  PCOUT(33) => R1IN_2_2_1_0(33),
  PCOUT(34) => UC_103_0,
  PCOUT(35) => UC_104_0,
  PCOUT(36) => UC_105_0,
  PCOUT(37) => UC_106_0,
  PCOUT(38) => UC_107_0,
  PCOUT(39) => UC_108_0,
  PCOUT(40) => UC_109_0,
  PCOUT(41) => UC_110_0,
  PCOUT(42) => UC_111_0,
  PCOUT(43) => UC_112_0,
  PCOUT(44) => UC_113_0,
  PCOUT(45) => UC_114_0,
  PCOUT(46) => UC_115_0,
  PCOUT(47) => UC_116_0);
\R1IN_4_3_ADD_1[26:0]\: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 1,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => B(51),
  A(1) => B(52),
  A(2) => B(53),
  A(3) => B(54),
  A(4) => B(55),
  A(5) => B(56),
  A(6) => B(57),
  A(7) => B(58),
  A(8) => B(59),
  A(9) => B(60),
  A(10) => NN_1,
  A(11) => NN_1,
  A(12) => NN_1,
  A(13) => NN_1,
  A(14) => NN_1,
  A(15) => NN_1,
  A(16) => NN_1,
  A(17) => NN_1,
  B(0) => A(17),
  B(1) => A(18),
  B(2) => A(19),
  B(3) => A(20),
  B(4) => A(21),
  B(5) => A(22),
  B(6) => A(23),
  B(7) => A(24),
  B(8) => A(25),
  B(9) => A(26),
  B(10) => A(27),
  B(11) => A(28),
  B(12) => A(29),
  B(13) => A(30),
  B(14) => A(31),
  B(15) => A(32),
  B(16) => A(33),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => R1IN_4_3_0(0),
  PCIN(1) => R1IN_4_3_0(1),
  PCIN(2) => R1IN_4_3_0(2),
  PCIN(3) => R1IN_4_3_0(3),
  PCIN(4) => R1IN_4_3_0(4),
  PCIN(5) => R1IN_4_3_0(5),
  PCIN(6) => R1IN_4_3_0(6),
  PCIN(7) => R1IN_4_3_0(7),
  PCIN(8) => R1IN_4_3_0(8),
  PCIN(9) => R1IN_4_3_0(9),
  PCIN(10) => R1IN_4_3_0(10),
  PCIN(11) => R1IN_4_3_0(11),
  PCIN(12) => R1IN_4_3_0(12),
  PCIN(13) => R1IN_4_3_0(13),
  PCIN(14) => R1IN_4_3_0(14),
  PCIN(15) => R1IN_4_3_0(15),
  PCIN(16) => R1IN_4_3_0(16),
  PCIN(17) => R1IN_4_3_1_0(17),
  PCIN(18) => R1IN_4_3_1_0(18),
  PCIN(19) => R1IN_4_3_1_0(19),
  PCIN(20) => R1IN_4_3_1_0(20),
  PCIN(21) => R1IN_4_3_1_0(21),
  PCIN(22) => R1IN_4_3_1_0(22),
  PCIN(23) => R1IN_4_3_1_0(23),
  PCIN(24) => R1IN_4_3_1_0(24),
  PCIN(25) => R1IN_4_3_1_0(25),
  PCIN(26) => R1IN_4_3_1_0(26),
  PCIN(27) => R1IN_4_3_1_0(27),
  PCIN(28) => R1IN_4_3_1_0(28),
  PCIN(29) => R1IN_4_3_1_0(29),
  PCIN(30) => R1IN_4_3_1_0(30),
  PCIN(31) => R1IN_4_3_1_0(31),
  PCIN(32) => R1IN_4_3_1_0(32),
  PCIN(33) => R1IN_4_3_1_0(33),
  PCIN(34) => UC_145_0,
  PCIN(35) => UC_146_0,
  PCIN(36) => UC_147_0,
  PCIN(37) => UC_148_0,
  PCIN(38) => UC_149_0,
  PCIN(39) => UC_150_0,
  PCIN(40) => UC_151_0,
  PCIN(41) => UC_152_0,
  PCIN(42) => UC_153_0,
  PCIN(43) => UC_154_0,
  PCIN(44) => UC_155_0,
  PCIN(45) => UC_156_0,
  PCIN(46) => UC_157_0,
  PCIN(47) => UC_158_0,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_2,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_2,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => CLK,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => EN,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_4_3_ADD_1_BCOUT(0),
  BCOUT(1) => R1IN_4_3_ADD_1_BCOUT(1),
  BCOUT(2) => R1IN_4_3_ADD_1_BCOUT(2),
  BCOUT(3) => R1IN_4_3_ADD_1_BCOUT(3),
  BCOUT(4) => R1IN_4_3_ADD_1_BCOUT(4),
  BCOUT(5) => R1IN_4_3_ADD_1_BCOUT(5),
  BCOUT(6) => R1IN_4_3_ADD_1_BCOUT(6),
  BCOUT(7) => R1IN_4_3_ADD_1_BCOUT(7),
  BCOUT(8) => R1IN_4_3_ADD_1_BCOUT(8),
  BCOUT(9) => R1IN_4_3_ADD_1_BCOUT(9),
  BCOUT(10) => R1IN_4_3_ADD_1_BCOUT(10),
  BCOUT(11) => R1IN_4_3_ADD_1_BCOUT(11),
  BCOUT(12) => R1IN_4_3_ADD_1_BCOUT(12),
  BCOUT(13) => R1IN_4_3_ADD_1_BCOUT(13),
  BCOUT(14) => R1IN_4_3_ADD_1_BCOUT(14),
  BCOUT(15) => R1IN_4_3_ADD_1_BCOUT(15),
  BCOUT(16) => R1IN_4_3_ADD_1_BCOUT(16),
  BCOUT(17) => R1IN_4_3_ADD_1_BCOUT(17),
  P(0) => R1IN_4_3F(17),
  P(1) => R1IN_4_3F(18),
  P(2) => R1IN_4_3F(19),
  P(3) => R1IN_4_3F(20),
  P(4) => R1IN_4_3F(21),
  P(5) => R1IN_4_3F(22),
  P(6) => R1IN_4_3F(23),
  P(7) => R1IN_4_3F(24),
  P(8) => R1IN_4_3F(25),
  P(9) => R1IN_4_3F(26),
  P(10) => R1IN_4_3F(27),
  P(11) => R1IN_4_3F(28),
  P(12) => R1IN_4_3F(29),
  P(13) => R1IN_4_3F(30),
  P(14) => R1IN_4_3F(31),
  P(15) => R1IN_4_3F(32),
  P(16) => R1IN_4_3F(33),
  P(17) => R1IN_4_3F(34),
  P(18) => R1IN_4_3F(35),
  P(19) => R1IN_4_3F(36),
  P(20) => R1IN_4_3F(37),
  P(21) => R1IN_4_3F(38),
  P(22) => R1IN_4_3F(39),
  P(23) => R1IN_4_3F(40),
  P(24) => R1IN_4_3F(41),
  P(25) => R1IN_4_3F(42),
  P(26) => R1IN_4_3F(43),
  P(27) => UC_82,
  P(28) => UC_83,
  P(29) => UC_84,
  P(30) => UC_85,
  P(31) => UC_86,
  P(32) => UC_87,
  P(33) => UC_88,
  P(34) => UC_89,
  P(35) => UC_90,
  P(36) => UC_91,
  P(37) => UC_92,
  P(38) => UC_93,
  P(39) => UC_94,
  P(40) => UC_95,
  P(41) => UC_96,
  P(42) => UC_97,
  P(43) => UC_98,
  P(44) => UC_99,
  P(45) => UC_100,
  P(46) => UC_101,
  P(47) => UC_102,
  PCOUT(0) => R1IN_4_3_ADD_1_PCOUT(0),
  PCOUT(1) => R1IN_4_3_ADD_1_PCOUT(1),
  PCOUT(2) => R1IN_4_3_ADD_1_PCOUT(2),
  PCOUT(3) => R1IN_4_3_ADD_1_PCOUT(3),
  PCOUT(4) => R1IN_4_3_ADD_1_PCOUT(4),
  PCOUT(5) => R1IN_4_3_ADD_1_PCOUT(5),
  PCOUT(6) => R1IN_4_3_ADD_1_PCOUT(6),
  PCOUT(7) => R1IN_4_3_ADD_1_PCOUT(7),
  PCOUT(8) => R1IN_4_3_ADD_1_PCOUT(8),
  PCOUT(9) => R1IN_4_3_ADD_1_PCOUT(9),
  PCOUT(10) => R1IN_4_3_ADD_1_PCOUT(10),
  PCOUT(11) => R1IN_4_3_ADD_1_PCOUT(11),
  PCOUT(12) => R1IN_4_3_ADD_1_PCOUT(12),
  PCOUT(13) => R1IN_4_3_ADD_1_PCOUT(13),
  PCOUT(14) => R1IN_4_3_ADD_1_PCOUT(14),
  PCOUT(15) => R1IN_4_3_ADD_1_PCOUT(15),
  PCOUT(16) => R1IN_4_3_ADD_1_PCOUT(16),
  PCOUT(17) => R1IN_4_3_ADD_1_PCOUT(17),
  PCOUT(18) => R1IN_4_3_ADD_1_PCOUT(18),
  PCOUT(19) => R1IN_4_3_ADD_1_PCOUT(19),
  PCOUT(20) => R1IN_4_3_ADD_1_PCOUT(20),
  PCOUT(21) => R1IN_4_3_ADD_1_PCOUT(21),
  PCOUT(22) => R1IN_4_3_ADD_1_PCOUT(22),
  PCOUT(23) => R1IN_4_3_ADD_1_PCOUT(23),
  PCOUT(24) => R1IN_4_3_ADD_1_PCOUT(24),
  PCOUT(25) => R1IN_4_3_ADD_1_PCOUT(25),
  PCOUT(26) => R1IN_4_3_ADD_1_PCOUT(26),
  PCOUT(27) => R1IN_4_3_ADD_1_PCOUT(27),
  PCOUT(28) => R1IN_4_3_ADD_1_PCOUT(28),
  PCOUT(29) => R1IN_4_3_ADD_1_PCOUT(29),
  PCOUT(30) => R1IN_4_3_ADD_1_PCOUT(30),
  PCOUT(31) => R1IN_4_3_ADD_1_PCOUT(31),
  PCOUT(32) => R1IN_4_3_ADD_1_PCOUT(32),
  PCOUT(33) => R1IN_4_3_ADD_1_PCOUT(33),
  PCOUT(34) => R1IN_4_3_ADD_1_PCOUT(34),
  PCOUT(35) => R1IN_4_3_ADD_1_PCOUT(35),
  PCOUT(36) => R1IN_4_3_ADD_1_PCOUT(36),
  PCOUT(37) => R1IN_4_3_ADD_1_PCOUT(37),
  PCOUT(38) => R1IN_4_3_ADD_1_PCOUT(38),
  PCOUT(39) => R1IN_4_3_ADD_1_PCOUT(39),
  PCOUT(40) => R1IN_4_3_ADD_1_PCOUT(40),
  PCOUT(41) => R1IN_4_3_ADD_1_PCOUT(41),
  PCOUT(42) => R1IN_4_3_ADD_1_PCOUT(42),
  PCOUT(43) => R1IN_4_3_ADD_1_PCOUT(43),
  PCOUT(44) => R1IN_4_3_ADD_1_PCOUT(44),
  PCOUT(45) => R1IN_4_3_ADD_1_PCOUT(45),
  PCOUT(46) => R1IN_4_3_ADD_1_PCOUT(46),
  PCOUT(47) => R1IN_4_3_ADD_1_PCOUT(47));
\R1IN_4_2_ADD_1[26:0]\: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 1,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => A(51),
  A(1) => A(52),
  A(2) => A(53),
  A(3) => A(54),
  A(4) => A(55),
  A(5) => A(56),
  A(6) => A(57),
  A(7) => A(58),
  A(8) => A(59),
  A(9) => A(60),
  A(10) => NN_1,
  A(11) => NN_1,
  A(12) => NN_1,
  A(13) => NN_1,
  A(14) => NN_1,
  A(15) => NN_1,
  A(16) => NN_1,
  A(17) => NN_1,
  B(0) => B(17),
  B(1) => B(18),
  B(2) => B(19),
  B(3) => B(20),
  B(4) => B(21),
  B(5) => B(22),
  B(6) => B(23),
  B(7) => B(24),
  B(8) => B(25),
  B(9) => B(26),
  B(10) => B(27),
  B(11) => B(28),
  B(12) => B(29),
  B(13) => B(30),
  B(14) => B(31),
  B(15) => B(32),
  B(16) => B(33),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => R1IN_4_2_0(0),
  PCIN(1) => R1IN_4_2_0(1),
  PCIN(2) => R1IN_4_2_0(2),
  PCIN(3) => R1IN_4_2_0(3),
  PCIN(4) => R1IN_4_2_0(4),
  PCIN(5) => R1IN_4_2_0(5),
  PCIN(6) => R1IN_4_2_0(6),
  PCIN(7) => R1IN_4_2_0(7),
  PCIN(8) => R1IN_4_2_0(8),
  PCIN(9) => R1IN_4_2_0(9),
  PCIN(10) => R1IN_4_2_0(10),
  PCIN(11) => R1IN_4_2_0(11),
  PCIN(12) => R1IN_4_2_0(12),
  PCIN(13) => R1IN_4_2_0(13),
  PCIN(14) => R1IN_4_2_0(14),
  PCIN(15) => R1IN_4_2_0(15),
  PCIN(16) => R1IN_4_2_0(16),
  PCIN(17) => R1IN_4_2_1_0(17),
  PCIN(18) => R1IN_4_2_1_0(18),
  PCIN(19) => R1IN_4_2_1_0(19),
  PCIN(20) => R1IN_4_2_1_0(20),
  PCIN(21) => R1IN_4_2_1_0(21),
  PCIN(22) => R1IN_4_2_1_0(22),
  PCIN(23) => R1IN_4_2_1_0(23),
  PCIN(24) => R1IN_4_2_1_0(24),
  PCIN(25) => R1IN_4_2_1_0(25),
  PCIN(26) => R1IN_4_2_1_0(26),
  PCIN(27) => R1IN_4_2_1_0(27),
  PCIN(28) => R1IN_4_2_1_0(28),
  PCIN(29) => R1IN_4_2_1_0(29),
  PCIN(30) => R1IN_4_2_1_0(30),
  PCIN(31) => R1IN_4_2_1_0(31),
  PCIN(32) => R1IN_4_2_1_0(32),
  PCIN(33) => R1IN_4_2_1_0(33),
  PCIN(34) => UC_131_0,
  PCIN(35) => UC_132_0,
  PCIN(36) => UC_133_0,
  PCIN(37) => UC_134_0,
  PCIN(38) => UC_135_0,
  PCIN(39) => UC_136_0,
  PCIN(40) => UC_137_0,
  PCIN(41) => UC_138_0,
  PCIN(42) => UC_139_0,
  PCIN(43) => UC_140_0,
  PCIN(44) => UC_141_0,
  PCIN(45) => UC_142_0,
  PCIN(46) => UC_143_0,
  PCIN(47) => UC_144_0,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_2,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_2,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => CLK,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => EN,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_4_2_ADD_1_BCOUT(0),
  BCOUT(1) => R1IN_4_2_ADD_1_BCOUT(1),
  BCOUT(2) => R1IN_4_2_ADD_1_BCOUT(2),
  BCOUT(3) => R1IN_4_2_ADD_1_BCOUT(3),
  BCOUT(4) => R1IN_4_2_ADD_1_BCOUT(4),
  BCOUT(5) => R1IN_4_2_ADD_1_BCOUT(5),
  BCOUT(6) => R1IN_4_2_ADD_1_BCOUT(6),
  BCOUT(7) => R1IN_4_2_ADD_1_BCOUT(7),
  BCOUT(8) => R1IN_4_2_ADD_1_BCOUT(8),
  BCOUT(9) => R1IN_4_2_ADD_1_BCOUT(9),
  BCOUT(10) => R1IN_4_2_ADD_1_BCOUT(10),
  BCOUT(11) => R1IN_4_2_ADD_1_BCOUT(11),
  BCOUT(12) => R1IN_4_2_ADD_1_BCOUT(12),
  BCOUT(13) => R1IN_4_2_ADD_1_BCOUT(13),
  BCOUT(14) => R1IN_4_2_ADD_1_BCOUT(14),
  BCOUT(15) => R1IN_4_2_ADD_1_BCOUT(15),
  BCOUT(16) => R1IN_4_2_ADD_1_BCOUT(16),
  BCOUT(17) => R1IN_4_2_ADD_1_BCOUT(17),
  P(0) => R1IN_4_2F(17),
  P(1) => R1IN_4_2F(18),
  P(2) => R1IN_4_2F(19),
  P(3) => R1IN_4_2F(20),
  P(4) => R1IN_4_2F(21),
  P(5) => R1IN_4_2F(22),
  P(6) => R1IN_4_2F(23),
  P(7) => R1IN_4_2F(24),
  P(8) => R1IN_4_2F(25),
  P(9) => R1IN_4_2F(26),
  P(10) => R1IN_4_2F(27),
  P(11) => R1IN_4_2F(28),
  P(12) => R1IN_4_2F(29),
  P(13) => R1IN_4_2F(30),
  P(14) => R1IN_4_2F(31),
  P(15) => R1IN_4_2F(32),
  P(16) => R1IN_4_2F(33),
  P(17) => R1IN_4_2F(34),
  P(18) => R1IN_4_2F(35),
  P(19) => R1IN_4_2F(36),
  P(20) => R1IN_4_2F(37),
  P(21) => R1IN_4_2F(38),
  P(22) => R1IN_4_2F(39),
  P(23) => R1IN_4_2F(40),
  P(24) => R1IN_4_2F(41),
  P(25) => R1IN_4_2F(42),
  P(26) => R1IN_4_2F(43),
  P(27) => UC_61,
  P(28) => UC_62,
  P(29) => UC_63,
  P(30) => UC_64,
  P(31) => UC_65,
  P(32) => UC_66,
  P(33) => UC_67,
  P(34) => UC_68,
  P(35) => UC_69,
  P(36) => UC_70,
  P(37) => UC_71,
  P(38) => UC_72,
  P(39) => UC_73,
  P(40) => UC_74,
  P(41) => UC_75,
  P(42) => UC_76,
  P(43) => UC_77,
  P(44) => UC_78,
  P(45) => UC_79,
  P(46) => UC_80,
  P(47) => UC_81,
  PCOUT(0) => R1IN_4_2_ADD_1_PCOUT(0),
  PCOUT(1) => R1IN_4_2_ADD_1_PCOUT(1),
  PCOUT(2) => R1IN_4_2_ADD_1_PCOUT(2),
  PCOUT(3) => R1IN_4_2_ADD_1_PCOUT(3),
  PCOUT(4) => R1IN_4_2_ADD_1_PCOUT(4),
  PCOUT(5) => R1IN_4_2_ADD_1_PCOUT(5),
  PCOUT(6) => R1IN_4_2_ADD_1_PCOUT(6),
  PCOUT(7) => R1IN_4_2_ADD_1_PCOUT(7),
  PCOUT(8) => R1IN_4_2_ADD_1_PCOUT(8),
  PCOUT(9) => R1IN_4_2_ADD_1_PCOUT(9),
  PCOUT(10) => R1IN_4_2_ADD_1_PCOUT(10),
  PCOUT(11) => R1IN_4_2_ADD_1_PCOUT(11),
  PCOUT(12) => R1IN_4_2_ADD_1_PCOUT(12),
  PCOUT(13) => R1IN_4_2_ADD_1_PCOUT(13),
  PCOUT(14) => R1IN_4_2_ADD_1_PCOUT(14),
  PCOUT(15) => R1IN_4_2_ADD_1_PCOUT(15),
  PCOUT(16) => R1IN_4_2_ADD_1_PCOUT(16),
  PCOUT(17) => R1IN_4_2_ADD_1_PCOUT(17),
  PCOUT(18) => R1IN_4_2_ADD_1_PCOUT(18),
  PCOUT(19) => R1IN_4_2_ADD_1_PCOUT(19),
  PCOUT(20) => R1IN_4_2_ADD_1_PCOUT(20),
  PCOUT(21) => R1IN_4_2_ADD_1_PCOUT(21),
  PCOUT(22) => R1IN_4_2_ADD_1_PCOUT(22),
  PCOUT(23) => R1IN_4_2_ADD_1_PCOUT(23),
  PCOUT(24) => R1IN_4_2_ADD_1_PCOUT(24),
  PCOUT(25) => R1IN_4_2_ADD_1_PCOUT(25),
  PCOUT(26) => R1IN_4_2_ADD_1_PCOUT(26),
  PCOUT(27) => R1IN_4_2_ADD_1_PCOUT(27),
  PCOUT(28) => R1IN_4_2_ADD_1_PCOUT(28),
  PCOUT(29) => R1IN_4_2_ADD_1_PCOUT(29),
  PCOUT(30) => R1IN_4_2_ADD_1_PCOUT(30),
  PCOUT(31) => R1IN_4_2_ADD_1_PCOUT(31),
  PCOUT(32) => R1IN_4_2_ADD_1_PCOUT(32),
  PCOUT(33) => R1IN_4_2_ADD_1_PCOUT(33),
  PCOUT(34) => R1IN_4_2_ADD_1_PCOUT(34),
  PCOUT(35) => R1IN_4_2_ADD_1_PCOUT(35),
  PCOUT(36) => R1IN_4_2_ADD_1_PCOUT(36),
  PCOUT(37) => R1IN_4_2_ADD_1_PCOUT(37),
  PCOUT(38) => R1IN_4_2_ADD_1_PCOUT(38),
  PCOUT(39) => R1IN_4_2_ADD_1_PCOUT(39),
  PCOUT(40) => R1IN_4_2_ADD_1_PCOUT(40),
  PCOUT(41) => R1IN_4_2_ADD_1_PCOUT(41),
  PCOUT(42) => R1IN_4_2_ADD_1_PCOUT(42),
  PCOUT(43) => R1IN_4_2_ADD_1_PCOUT(43),
  PCOUT(44) => R1IN_4_2_ADD_1_PCOUT(44),
  PCOUT(45) => R1IN_4_2_ADD_1_PCOUT(45),
  PCOUT(46) => R1IN_4_2_ADD_1_PCOUT(46),
  PCOUT(47) => R1IN_4_2_ADD_1_PCOUT(47));
\R1IN_3_2_ADD_1[26:0]\: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 1,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => B(51),
  A(1) => B(52),
  A(2) => B(53),
  A(3) => B(54),
  A(4) => B(55),
  A(5) => B(56),
  A(6) => B(57),
  A(7) => B(58),
  A(8) => B(59),
  A(9) => B(60),
  A(10) => NN_1,
  A(11) => NN_1,
  A(12) => NN_1,
  A(13) => NN_1,
  A(14) => NN_1,
  A(15) => NN_1,
  A(16) => NN_1,
  A(17) => NN_1,
  B(0) => A(0),
  B(1) => A(1),
  B(2) => A(2),
  B(3) => A(3),
  B(4) => A(4),
  B(5) => A(5),
  B(6) => A(6),
  B(7) => A(7),
  B(8) => A(8),
  B(9) => A(9),
  B(10) => A(10),
  B(11) => A(11),
  B(12) => A(12),
  B(13) => A(13),
  B(14) => A(14),
  B(15) => A(15),
  B(16) => A(16),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => R1IN_3_2_0(0),
  PCIN(1) => R1IN_3_2_0(1),
  PCIN(2) => R1IN_3_2_0(2),
  PCIN(3) => R1IN_3_2_0(3),
  PCIN(4) => R1IN_3_2_0(4),
  PCIN(5) => R1IN_3_2_0(5),
  PCIN(6) => R1IN_3_2_0(6),
  PCIN(7) => R1IN_3_2_0(7),
  PCIN(8) => R1IN_3_2_0(8),
  PCIN(9) => R1IN_3_2_0(9),
  PCIN(10) => R1IN_3_2_0(10),
  PCIN(11) => R1IN_3_2_0(11),
  PCIN(12) => R1IN_3_2_0(12),
  PCIN(13) => R1IN_3_2_0(13),
  PCIN(14) => R1IN_3_2_0(14),
  PCIN(15) => R1IN_3_2_0(15),
  PCIN(16) => R1IN_3_2_0(16),
  PCIN(17) => R1IN_3_2_1_0(17),
  PCIN(18) => R1IN_3_2_1_0(18),
  PCIN(19) => R1IN_3_2_1_0(19),
  PCIN(20) => R1IN_3_2_1_0(20),
  PCIN(21) => R1IN_3_2_1_0(21),
  PCIN(22) => R1IN_3_2_1_0(22),
  PCIN(23) => R1IN_3_2_1_0(23),
  PCIN(24) => R1IN_3_2_1_0(24),
  PCIN(25) => R1IN_3_2_1_0(25),
  PCIN(26) => R1IN_3_2_1_0(26),
  PCIN(27) => R1IN_3_2_1_0(27),
  PCIN(28) => R1IN_3_2_1_0(28),
  PCIN(29) => R1IN_3_2_1_0(29),
  PCIN(30) => R1IN_3_2_1_0(30),
  PCIN(31) => R1IN_3_2_1_0(31),
  PCIN(32) => R1IN_3_2_1_0(32),
  PCIN(33) => R1IN_3_2_1_0(33),
  PCIN(34) => UC_117_0,
  PCIN(35) => UC_118_0,
  PCIN(36) => UC_119_0,
  PCIN(37) => UC_120_0,
  PCIN(38) => UC_121_0,
  PCIN(39) => UC_122_0,
  PCIN(40) => UC_123_0,
  PCIN(41) => UC_124_0,
  PCIN(42) => UC_125_0,
  PCIN(43) => UC_126_0,
  PCIN(44) => UC_127_0,
  PCIN(45) => UC_128_0,
  PCIN(46) => UC_129_0,
  PCIN(47) => UC_130_0,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_2,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_2,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => CLK,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => EN,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_3_2_ADD_1_BCOUT(0),
  BCOUT(1) => R1IN_3_2_ADD_1_BCOUT(1),
  BCOUT(2) => R1IN_3_2_ADD_1_BCOUT(2),
  BCOUT(3) => R1IN_3_2_ADD_1_BCOUT(3),
  BCOUT(4) => R1IN_3_2_ADD_1_BCOUT(4),
  BCOUT(5) => R1IN_3_2_ADD_1_BCOUT(5),
  BCOUT(6) => R1IN_3_2_ADD_1_BCOUT(6),
  BCOUT(7) => R1IN_3_2_ADD_1_BCOUT(7),
  BCOUT(8) => R1IN_3_2_ADD_1_BCOUT(8),
  BCOUT(9) => R1IN_3_2_ADD_1_BCOUT(9),
  BCOUT(10) => R1IN_3_2_ADD_1_BCOUT(10),
  BCOUT(11) => R1IN_3_2_ADD_1_BCOUT(11),
  BCOUT(12) => R1IN_3_2_ADD_1_BCOUT(12),
  BCOUT(13) => R1IN_3_2_ADD_1_BCOUT(13),
  BCOUT(14) => R1IN_3_2_ADD_1_BCOUT(14),
  BCOUT(15) => R1IN_3_2_ADD_1_BCOUT(15),
  BCOUT(16) => R1IN_3_2_ADD_1_BCOUT(16),
  BCOUT(17) => R1IN_3_2_ADD_1_BCOUT(17),
  P(0) => R1IN_3_2F(17),
  P(1) => R1IN_3_2F(18),
  P(2) => R1IN_3_2F(19),
  P(3) => R1IN_3_2F(20),
  P(4) => R1IN_3_2F(21),
  P(5) => R1IN_3_2F(22),
  P(6) => R1IN_3_2F(23),
  P(7) => R1IN_3_2F(24),
  P(8) => R1IN_3_2F(25),
  P(9) => R1IN_3_2F(26),
  P(10) => R1IN_3_2F(27),
  P(11) => R1IN_3_2F(28),
  P(12) => R1IN_3_2F(29),
  P(13) => R1IN_3_2F(30),
  P(14) => R1IN_3_2F(31),
  P(15) => R1IN_3_2F(32),
  P(16) => R1IN_3_2F(33),
  P(17) => R1IN_3_2F(34),
  P(18) => R1IN_3_2F(35),
  P(19) => R1IN_3_2F(36),
  P(20) => R1IN_3_2F(37),
  P(21) => R1IN_3_2F(38),
  P(22) => R1IN_3_2F(39),
  P(23) => R1IN_3_2F(40),
  P(24) => R1IN_3_2F(41),
  P(25) => R1IN_3_2F(42),
  P(26) => R1IN_3_2F(43),
  P(27) => UC_40,
  P(28) => UC_41,
  P(29) => UC_42,
  P(30) => UC_43,
  P(31) => UC_44,
  P(32) => UC_45,
  P(33) => UC_46,
  P(34) => UC_47,
  P(35) => UC_48,
  P(36) => UC_49,
  P(37) => UC_50,
  P(38) => UC_51,
  P(39) => UC_52,
  P(40) => UC_53,
  P(41) => UC_54,
  P(42) => UC_55,
  P(43) => UC_56,
  P(44) => UC_57,
  P(45) => UC_58,
  P(46) => UC_59,
  P(47) => UC_60,
  PCOUT(0) => R1IN_3_2_ADD_1_PCOUT(0),
  PCOUT(1) => R1IN_3_2_ADD_1_PCOUT(1),
  PCOUT(2) => R1IN_3_2_ADD_1_PCOUT(2),
  PCOUT(3) => R1IN_3_2_ADD_1_PCOUT(3),
  PCOUT(4) => R1IN_3_2_ADD_1_PCOUT(4),
  PCOUT(5) => R1IN_3_2_ADD_1_PCOUT(5),
  PCOUT(6) => R1IN_3_2_ADD_1_PCOUT(6),
  PCOUT(7) => R1IN_3_2_ADD_1_PCOUT(7),
  PCOUT(8) => R1IN_3_2_ADD_1_PCOUT(8),
  PCOUT(9) => R1IN_3_2_ADD_1_PCOUT(9),
  PCOUT(10) => R1IN_3_2_ADD_1_PCOUT(10),
  PCOUT(11) => R1IN_3_2_ADD_1_PCOUT(11),
  PCOUT(12) => R1IN_3_2_ADD_1_PCOUT(12),
  PCOUT(13) => R1IN_3_2_ADD_1_PCOUT(13),
  PCOUT(14) => R1IN_3_2_ADD_1_PCOUT(14),
  PCOUT(15) => R1IN_3_2_ADD_1_PCOUT(15),
  PCOUT(16) => R1IN_3_2_ADD_1_PCOUT(16),
  PCOUT(17) => R1IN_3_2_ADD_1_PCOUT(17),
  PCOUT(18) => R1IN_3_2_ADD_1_PCOUT(18),
  PCOUT(19) => R1IN_3_2_ADD_1_PCOUT(19),
  PCOUT(20) => R1IN_3_2_ADD_1_PCOUT(20),
  PCOUT(21) => R1IN_3_2_ADD_1_PCOUT(21),
  PCOUT(22) => R1IN_3_2_ADD_1_PCOUT(22),
  PCOUT(23) => R1IN_3_2_ADD_1_PCOUT(23),
  PCOUT(24) => R1IN_3_2_ADD_1_PCOUT(24),
  PCOUT(25) => R1IN_3_2_ADD_1_PCOUT(25),
  PCOUT(26) => R1IN_3_2_ADD_1_PCOUT(26),
  PCOUT(27) => R1IN_3_2_ADD_1_PCOUT(27),
  PCOUT(28) => R1IN_3_2_ADD_1_PCOUT(28),
  PCOUT(29) => R1IN_3_2_ADD_1_PCOUT(29),
  PCOUT(30) => R1IN_3_2_ADD_1_PCOUT(30),
  PCOUT(31) => R1IN_3_2_ADD_1_PCOUT(31),
  PCOUT(32) => R1IN_3_2_ADD_1_PCOUT(32),
  PCOUT(33) => R1IN_3_2_ADD_1_PCOUT(33),
  PCOUT(34) => R1IN_3_2_ADD_1_PCOUT(34),
  PCOUT(35) => R1IN_3_2_ADD_1_PCOUT(35),
  PCOUT(36) => R1IN_3_2_ADD_1_PCOUT(36),
  PCOUT(37) => R1IN_3_2_ADD_1_PCOUT(37),
  PCOUT(38) => R1IN_3_2_ADD_1_PCOUT(38),
  PCOUT(39) => R1IN_3_2_ADD_1_PCOUT(39),
  PCOUT(40) => R1IN_3_2_ADD_1_PCOUT(40),
  PCOUT(41) => R1IN_3_2_ADD_1_PCOUT(41),
  PCOUT(42) => R1IN_3_2_ADD_1_PCOUT(42),
  PCOUT(43) => R1IN_3_2_ADD_1_PCOUT(43),
  PCOUT(44) => R1IN_3_2_ADD_1_PCOUT(44),
  PCOUT(45) => R1IN_3_2_ADD_1_PCOUT(45),
  PCOUT(46) => R1IN_3_2_ADD_1_PCOUT(46),
  PCOUT(47) => R1IN_3_2_ADD_1_PCOUT(47));
\R1IN_2_2_ADD_1[26:0]\: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 1,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => A(51),
  A(1) => A(52),
  A(2) => A(53),
  A(3) => A(54),
  A(4) => A(55),
  A(5) => A(56),
  A(6) => A(57),
  A(7) => A(58),
  A(8) => A(59),
  A(9) => A(60),
  A(10) => NN_1,
  A(11) => NN_1,
  A(12) => NN_1,
  A(13) => NN_1,
  A(14) => NN_1,
  A(15) => NN_1,
  A(16) => NN_1,
  A(17) => NN_1,
  B(0) => B(0),
  B(1) => B(1),
  B(2) => B(2),
  B(3) => B(3),
  B(4) => B(4),
  B(5) => B(5),
  B(6) => B(6),
  B(7) => B(7),
  B(8) => B(8),
  B(9) => B(9),
  B(10) => B(10),
  B(11) => B(11),
  B(12) => B(12),
  B(13) => B(13),
  B(14) => B(14),
  B(15) => B(15),
  B(16) => B(16),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => R1IN_2_2_0(0),
  PCIN(1) => R1IN_2_2_0(1),
  PCIN(2) => R1IN_2_2_0(2),
  PCIN(3) => R1IN_2_2_0(3),
  PCIN(4) => R1IN_2_2_0(4),
  PCIN(5) => R1IN_2_2_0(5),
  PCIN(6) => R1IN_2_2_0(6),
  PCIN(7) => R1IN_2_2_0(7),
  PCIN(8) => R1IN_2_2_0(8),
  PCIN(9) => R1IN_2_2_0(9),
  PCIN(10) => R1IN_2_2_0(10),
  PCIN(11) => R1IN_2_2_0(11),
  PCIN(12) => R1IN_2_2_0(12),
  PCIN(13) => R1IN_2_2_0(13),
  PCIN(14) => R1IN_2_2_0(14),
  PCIN(15) => R1IN_2_2_0(15),
  PCIN(16) => R1IN_2_2_0(16),
  PCIN(17) => R1IN_2_2_1_0(17),
  PCIN(18) => R1IN_2_2_1_0(18),
  PCIN(19) => R1IN_2_2_1_0(19),
  PCIN(20) => R1IN_2_2_1_0(20),
  PCIN(21) => R1IN_2_2_1_0(21),
  PCIN(22) => R1IN_2_2_1_0(22),
  PCIN(23) => R1IN_2_2_1_0(23),
  PCIN(24) => R1IN_2_2_1_0(24),
  PCIN(25) => R1IN_2_2_1_0(25),
  PCIN(26) => R1IN_2_2_1_0(26),
  PCIN(27) => R1IN_2_2_1_0(27),
  PCIN(28) => R1IN_2_2_1_0(28),
  PCIN(29) => R1IN_2_2_1_0(29),
  PCIN(30) => R1IN_2_2_1_0(30),
  PCIN(31) => R1IN_2_2_1_0(31),
  PCIN(32) => R1IN_2_2_1_0(32),
  PCIN(33) => R1IN_2_2_1_0(33),
  PCIN(34) => UC_103_0,
  PCIN(35) => UC_104_0,
  PCIN(36) => UC_105_0,
  PCIN(37) => UC_106_0,
  PCIN(38) => UC_107_0,
  PCIN(39) => UC_108_0,
  PCIN(40) => UC_109_0,
  PCIN(41) => UC_110_0,
  PCIN(42) => UC_111_0,
  PCIN(43) => UC_112_0,
  PCIN(44) => UC_113_0,
  PCIN(45) => UC_114_0,
  PCIN(46) => UC_115_0,
  PCIN(47) => UC_116_0,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_2,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_2,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => CLK,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => EN,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => B_0(0),
  BCOUT(1) => B_0(1),
  BCOUT(2) => B_0(2),
  BCOUT(3) => B_0(3),
  BCOUT(4) => B_0(4),
  BCOUT(5) => B_0(5),
  BCOUT(6) => B_0(6),
  BCOUT(7) => B_0(7),
  BCOUT(8) => B_0(8),
  BCOUT(9) => B_0(9),
  BCOUT(10) => B_0(10),
  BCOUT(11) => B_0(11),
  BCOUT(12) => B_0(12),
  BCOUT(13) => B_0(13),
  BCOUT(14) => B_0(14),
  BCOUT(15) => B_0(15),
  BCOUT(16) => B_0(16),
  BCOUT(17) => GND_0,
  P(0) => R1IN_2_2F(17),
  P(1) => R1IN_2_2F(18),
  P(2) => R1IN_2_2F(19),
  P(3) => R1IN_2_2F(20),
  P(4) => R1IN_2_2F(21),
  P(5) => R1IN_2_2F(22),
  P(6) => R1IN_2_2F(23),
  P(7) => R1IN_2_2F(24),
  P(8) => R1IN_2_2F(25),
  P(9) => R1IN_2_2F(26),
  P(10) => R1IN_2_2F(27),
  P(11) => R1IN_2_2F(28),
  P(12) => R1IN_2_2F(29),
  P(13) => R1IN_2_2F(30),
  P(14) => R1IN_2_2F(31),
  P(15) => R1IN_2_2F(32),
  P(16) => R1IN_2_2F(33),
  P(17) => R1IN_2_2F(34),
  P(18) => R1IN_2_2F(35),
  P(19) => R1IN_2_2F(36),
  P(20) => R1IN_2_2F(37),
  P(21) => R1IN_2_2F(38),
  P(22) => R1IN_2_2F(39),
  P(23) => R1IN_2_2F(40),
  P(24) => R1IN_2_2F(41),
  P(25) => R1IN_2_2F(42),
  P(26) => R1IN_2_2F(43),
  P(27) => UC_19,
  P(28) => UC_20,
  P(29) => UC_21,
  P(30) => UC_22,
  P(31) => UC_23,
  P(32) => UC_24,
  P(33) => UC_25,
  P(34) => UC_26,
  P(35) => UC_27,
  P(36) => UC_28,
  P(37) => UC_29,
  P(38) => UC_30,
  P(39) => UC_31,
  P(40) => UC_32,
  P(41) => UC_33,
  P(42) => UC_34,
  P(43) => UC_35,
  P(44) => UC_36,
  P(45) => UC_37,
  P(46) => UC_38,
  P(47) => UC_39,
  PCOUT(0) => R1IN_2_2_ADD_1_PCOUT(0),
  PCOUT(1) => R1IN_2_2_ADD_1_PCOUT(1),
  PCOUT(2) => R1IN_2_2_ADD_1_PCOUT(2),
  PCOUT(3) => R1IN_2_2_ADD_1_PCOUT(3),
  PCOUT(4) => R1IN_2_2_ADD_1_PCOUT(4),
  PCOUT(5) => R1IN_2_2_ADD_1_PCOUT(5),
  PCOUT(6) => R1IN_2_2_ADD_1_PCOUT(6),
  PCOUT(7) => R1IN_2_2_ADD_1_PCOUT(7),
  PCOUT(8) => R1IN_2_2_ADD_1_PCOUT(8),
  PCOUT(9) => R1IN_2_2_ADD_1_PCOUT(9),
  PCOUT(10) => R1IN_2_2_ADD_1_PCOUT(10),
  PCOUT(11) => R1IN_2_2_ADD_1_PCOUT(11),
  PCOUT(12) => R1IN_2_2_ADD_1_PCOUT(12),
  PCOUT(13) => R1IN_2_2_ADD_1_PCOUT(13),
  PCOUT(14) => R1IN_2_2_ADD_1_PCOUT(14),
  PCOUT(15) => R1IN_2_2_ADD_1_PCOUT(15),
  PCOUT(16) => R1IN_2_2_ADD_1_PCOUT(16),
  PCOUT(17) => R1IN_2_2_ADD_1_PCOUT(17),
  PCOUT(18) => R1IN_2_2_ADD_1_PCOUT(18),
  PCOUT(19) => R1IN_2_2_ADD_1_PCOUT(19),
  PCOUT(20) => R1IN_2_2_ADD_1_PCOUT(20),
  PCOUT(21) => R1IN_2_2_ADD_1_PCOUT(21),
  PCOUT(22) => R1IN_2_2_ADD_1_PCOUT(22),
  PCOUT(23) => R1IN_2_2_ADD_1_PCOUT(23),
  PCOUT(24) => R1IN_2_2_ADD_1_PCOUT(24),
  PCOUT(25) => R1IN_2_2_ADD_1_PCOUT(25),
  PCOUT(26) => R1IN_2_2_ADD_1_PCOUT(26),
  PCOUT(27) => R1IN_2_2_ADD_1_PCOUT(27),
  PCOUT(28) => R1IN_2_2_ADD_1_PCOUT(28),
  PCOUT(29) => R1IN_2_2_ADD_1_PCOUT(29),
  PCOUT(30) => R1IN_2_2_ADD_1_PCOUT(30),
  PCOUT(31) => R1IN_2_2_ADD_1_PCOUT(31),
  PCOUT(32) => R1IN_2_2_ADD_1_PCOUT(32),
  PCOUT(33) => R1IN_2_2_ADD_1_PCOUT(33),
  PCOUT(34) => R1IN_2_2_ADD_1_PCOUT(34),
  PCOUT(35) => R1IN_2_2_ADD_1_PCOUT(35),
  PCOUT(36) => R1IN_2_2_ADD_1_PCOUT(36),
  PCOUT(37) => R1IN_2_2_ADD_1_PCOUT(37),
  PCOUT(38) => R1IN_2_2_ADD_1_PCOUT(38),
  PCOUT(39) => R1IN_2_2_ADD_1_PCOUT(39),
  PCOUT(40) => R1IN_2_2_ADD_1_PCOUT(40),
  PCOUT(41) => R1IN_2_2_ADD_1_PCOUT(41),
  PCOUT(42) => R1IN_2_2_ADD_1_PCOUT(42),
  PCOUT(43) => R1IN_2_2_ADD_1_PCOUT(43),
  PCOUT(44) => R1IN_2_2_ADD_1_PCOUT(44),
  PCOUT(45) => R1IN_2_2_ADD_1_PCOUT(45),
  PCOUT(46) => R1IN_2_2_ADD_1_PCOUT(46),
  PCOUT(47) => R1IN_2_2_ADD_1_PCOUT(47));
\R1IN_4_4_ADD_1[27:0]\: DSP48 
generic map(
  AREG => 0,
  BREG => 0,
  CREG => 0,
  PREG => 1,
  MREG => 0,
  SUBTRACTREG => 0,
  OPMODEREG => 0,
  CARRYINSELREG => 0,
  CARRYINREG => 0,
  B_INPUT => "DIRECT",
  LEGACY_MODE => "MULT18X18"
)
port map (
  A(0) => B(51),
  A(1) => B(52),
  A(2) => B(53),
  A(3) => B(54),
  A(4) => B(55),
  A(5) => B(56),
  A(6) => B(57),
  A(7) => B(58),
  A(8) => B(59),
  A(9) => B(60),
  A(10) => NN_1,
  A(11) => NN_1,
  A(12) => NN_1,
  A(13) => NN_1,
  A(14) => NN_1,
  A(15) => NN_1,
  A(16) => NN_1,
  A(17) => NN_1,
  B(0) => A(34),
  B(1) => A(35),
  B(2) => A(36),
  B(3) => A(37),
  B(4) => A(38),
  B(5) => A(39),
  B(6) => A(40),
  B(7) => A(41),
  B(8) => A(42),
  B(9) => A(43),
  B(10) => A(44),
  B(11) => A(45),
  B(12) => A(46),
  B(13) => A(47),
  B(14) => A(48),
  B(15) => A(49),
  B(16) => A(50),
  B(17) => NN_1,
  C(0) => NN_1,
  C(1) => NN_1,
  C(2) => NN_1,
  C(3) => NN_1,
  C(4) => NN_1,
  C(5) => NN_1,
  C(6) => NN_1,
  C(7) => NN_1,
  C(8) => NN_1,
  C(9) => NN_1,
  C(10) => NN_1,
  C(11) => NN_1,
  C(12) => NN_1,
  C(13) => NN_1,
  C(14) => NN_1,
  C(15) => NN_1,
  C(16) => NN_1,
  C(17) => NN_1,
  C(18) => NN_1,
  C(19) => NN_1,
  C(20) => NN_1,
  C(21) => NN_1,
  C(22) => NN_1,
  C(23) => NN_1,
  C(24) => NN_1,
  C(25) => NN_1,
  C(26) => NN_1,
  C(27) => NN_1,
  C(28) => NN_1,
  C(29) => NN_1,
  C(30) => NN_1,
  C(31) => NN_1,
  C(32) => NN_1,
  C(33) => NN_1,
  C(34) => NN_1,
  C(35) => NN_1,
  C(36) => NN_1,
  C(37) => NN_1,
  C(38) => NN_1,
  C(39) => NN_1,
  C(40) => NN_1,
  C(41) => NN_1,
  C(42) => NN_1,
  C(43) => NN_1,
  C(44) => NN_1,
  C(45) => NN_1,
  C(46) => NN_1,
  C(47) => NN_1,
  BCIN(0) => NN_1,
  BCIN(1) => NN_1,
  BCIN(2) => NN_1,
  BCIN(3) => NN_1,
  BCIN(4) => NN_1,
  BCIN(5) => NN_1,
  BCIN(6) => NN_1,
  BCIN(7) => NN_1,
  BCIN(8) => NN_1,
  BCIN(9) => NN_1,
  BCIN(10) => NN_1,
  BCIN(11) => NN_1,
  BCIN(12) => NN_1,
  BCIN(13) => NN_1,
  BCIN(14) => NN_1,
  BCIN(15) => NN_1,
  BCIN(16) => NN_1,
  BCIN(17) => NN_1,
  PCIN(0) => R1IN_4_4_2_0(0),
  PCIN(1) => R1IN_4_4_2_0(1),
  PCIN(2) => R1IN_4_4_2_0(2),
  PCIN(3) => R1IN_4_4_2_0(3),
  PCIN(4) => R1IN_4_4_2_0(4),
  PCIN(5) => R1IN_4_4_2_0(5),
  PCIN(6) => R1IN_4_4_2_0(6),
  PCIN(7) => R1IN_4_4_2_0(7),
  PCIN(8) => R1IN_4_4_2_0(8),
  PCIN(9) => R1IN_4_4_2_0(9),
  PCIN(10) => R1IN_4_4_2_0(10),
  PCIN(11) => R1IN_4_4_2_0(11),
  PCIN(12) => R1IN_4_4_2_0(12),
  PCIN(13) => R1IN_4_4_2_0(13),
  PCIN(14) => R1IN_4_4_2_0(14),
  PCIN(15) => R1IN_4_4_2_0(15),
  PCIN(16) => R1IN_4_4_2_0(16),
  PCIN(17) => R1IN_4_4_2_0(17),
  PCIN(18) => R1IN_4_4_2_0(18),
  PCIN(19) => R1IN_4_4_2_0(19),
  PCIN(20) => R1IN_4_4_2_0(20),
  PCIN(21) => R1IN_4_4_2_0(21),
  PCIN(22) => R1IN_4_4_2_0(22),
  PCIN(23) => R1IN_4_4_2_0(23),
  PCIN(24) => R1IN_4_4_2_0(24),
  PCIN(25) => R1IN_4_4_2_0(25),
  PCIN(26) => R1IN_4_4_2_0(26),
  PCIN(27) => UC_229_0,
  PCIN(28) => UC_230_0,
  PCIN(29) => UC_231_0,
  PCIN(30) => UC_232_0,
  PCIN(31) => UC_233_0,
  PCIN(32) => UC_234_0,
  PCIN(33) => UC_235_0,
  PCIN(34) => UC_236_0,
  PCIN(35) => UC_237_0,
  PCIN(36) => UC_238_0,
  PCIN(37) => UC_239_0,
  PCIN(38) => UC_240_0,
  PCIN(39) => UC_241_0,
  PCIN(40) => UC_242_0,
  PCIN(41) => UC_243_0,
  PCIN(42) => UC_244_0,
  PCIN(43) => UC_245_0,
  PCIN(44) => UC_246_0,
  PCIN(45) => UC_247_0,
  PCIN(46) => UC_248_0,
  PCIN(47) => UC_249_0,
  OPMODE(0) => NN_2,
  OPMODE(1) => NN_1,
  OPMODE(2) => NN_2,
  OPMODE(3) => NN_1,
  OPMODE(4) => NN_2,
  OPMODE(5) => NN_1,
  OPMODE(6) => NN_1,
  SUBTRACT => NN_1,
  CARRYIN => NN_1,
  CARRYINSEL(0) => NN_1,
  CARRYINSEL(1) => NN_1,
  CLK => CLK,
  CEA => NN_1,
  CEB => NN_1,
  CEC => NN_1,
  CEP => EN,
  CEM => NN_1,
  CECARRYIN => NN_1,
  CECTRL => NN_1,
  CECINSUB => NN_1,
  RSTA => NN_1,
  RSTB => NN_1,
  RSTC => NN_1,
  RSTP => NN_1,
  RSTM => NN_1,
  RSTCTRL => NN_1,
  RSTCARRYIN => NN_1,
  BCOUT(0) => R1IN_4_4_ADD_1_BCOUT(0),
  BCOUT(1) => R1IN_4_4_ADD_1_BCOUT(1),
  BCOUT(2) => R1IN_4_4_ADD_1_BCOUT(2),
  BCOUT(3) => R1IN_4_4_ADD_1_BCOUT(3),
  BCOUT(4) => R1IN_4_4_ADD_1_BCOUT(4),
  BCOUT(5) => R1IN_4_4_ADD_1_BCOUT(5),
  BCOUT(6) => R1IN_4_4_ADD_1_BCOUT(6),
  BCOUT(7) => R1IN_4_4_ADD_1_BCOUT(7),
  BCOUT(8) => R1IN_4_4_ADD_1_BCOUT(8),
  BCOUT(9) => R1IN_4_4_ADD_1_BCOUT(9),
  BCOUT(10) => R1IN_4_4_ADD_1_BCOUT(10),
  BCOUT(11) => R1IN_4_4_ADD_1_BCOUT(11),
  BCOUT(12) => R1IN_4_4_ADD_1_BCOUT(12),
  BCOUT(13) => R1IN_4_4_ADD_1_BCOUT(13),
  BCOUT(14) => R1IN_4_4_ADD_1_BCOUT(14),
  BCOUT(15) => R1IN_4_4_ADD_1_BCOUT(15),
  BCOUT(16) => R1IN_4_4_ADD_1_BCOUT(16),
  BCOUT(17) => R1IN_4_4_ADD_1_BCOUT(17),
  P(0) => R1IN_4_4_ADD_1F(0),
  P(1) => R1IN_4_4_ADD_1F(1),
  P(2) => R1IN_4_4_ADD_1F(2),
  P(3) => R1IN_4_4_ADD_1F(3),
  P(4) => R1IN_4_4_ADD_1F(4),
  P(5) => R1IN_4_4_ADD_1F(5),
  P(6) => R1IN_4_4_ADD_1F(6),
  P(7) => R1IN_4_4_ADD_1F(7),
  P(8) => R1IN_4_4_ADD_1F(8),
  P(9) => R1IN_4_4_ADD_1F(9),
  P(10) => R1IN_4_4_ADD_1F(10),
  P(11) => R1IN_4_4_ADD_1F(11),
  P(12) => R1IN_4_4_ADD_1F(12),
  P(13) => R1IN_4_4_ADD_1F(13),
  P(14) => R1IN_4_4_ADD_1F(14),
  P(15) => R1IN_4_4_ADD_1F(15),
  P(16) => R1IN_4_4_ADD_1F(16),
  P(17) => R1IN_4_4_ADD_1F(17),
  P(18) => R1IN_4_4_ADD_1F(18),
  P(19) => R1IN_4_4_ADD_1F(19),
  P(20) => R1IN_4_4_ADD_1F(20),
  P(21) => R1IN_4_4_ADD_1F(21),
  P(22) => R1IN_4_4_ADD_1F(22),
  P(23) => R1IN_4_4_ADD_1F(23),
  P(24) => R1IN_4_4_ADD_1F(24),
  P(25) => R1IN_4_4_ADD_1F(25),
  P(26) => R1IN_4_4_ADD_1F(26),
  P(27) => R1IN_4_4_ADD_1F(27),
  P(28) => UC,
  P(29) => UC_0,
  P(30) => UC_1,
  P(31) => UC_2,
  P(32) => UC_3,
  P(33) => UC_4,
  P(34) => UC_5,
  P(35) => UC_6,
  P(36) => UC_7,
  P(37) => UC_8,
  P(38) => UC_9,
  P(39) => UC_10,
  P(40) => UC_11,
  P(41) => UC_12,
  P(42) => UC_13,
  P(43) => UC_14,
  P(44) => UC_15,
  P(45) => UC_16,
  P(46) => UC_17,
  P(47) => UC_18,
  PCOUT(0) => R1IN_4_4_ADD_1_PCOUT(0),
  PCOUT(1) => R1IN_4_4_ADD_1_PCOUT(1),
  PCOUT(2) => R1IN_4_4_ADD_1_PCOUT(2),
  PCOUT(3) => R1IN_4_4_ADD_1_PCOUT(3),
  PCOUT(4) => R1IN_4_4_ADD_1_PCOUT(4),
  PCOUT(5) => R1IN_4_4_ADD_1_PCOUT(5),
  PCOUT(6) => R1IN_4_4_ADD_1_PCOUT(6),
  PCOUT(7) => R1IN_4_4_ADD_1_PCOUT(7),
  PCOUT(8) => R1IN_4_4_ADD_1_PCOUT(8),
  PCOUT(9) => R1IN_4_4_ADD_1_PCOUT(9),
  PCOUT(10) => R1IN_4_4_ADD_1_PCOUT(10),
  PCOUT(11) => R1IN_4_4_ADD_1_PCOUT(11),
  PCOUT(12) => R1IN_4_4_ADD_1_PCOUT(12),
  PCOUT(13) => R1IN_4_4_ADD_1_PCOUT(13),
  PCOUT(14) => R1IN_4_4_ADD_1_PCOUT(14),
  PCOUT(15) => R1IN_4_4_ADD_1_PCOUT(15),
  PCOUT(16) => R1IN_4_4_ADD_1_PCOUT(16),
  PCOUT(17) => R1IN_4_4_ADD_1_PCOUT(17),
  PCOUT(18) => R1IN_4_4_ADD_1_PCOUT(18),
  PCOUT(19) => R1IN_4_4_ADD_1_PCOUT(19),
  PCOUT(20) => R1IN_4_4_ADD_1_PCOUT(20),
  PCOUT(21) => R1IN_4_4_ADD_1_PCOUT(21),
  PCOUT(22) => R1IN_4_4_ADD_1_PCOUT(22),
  PCOUT(23) => R1IN_4_4_ADD_1_PCOUT(23),
  PCOUT(24) => R1IN_4_4_ADD_1_PCOUT(24),
  PCOUT(25) => R1IN_4_4_ADD_1_PCOUT(25),
  PCOUT(26) => R1IN_4_4_ADD_1_PCOUT(26),
  PCOUT(27) => R1IN_4_4_ADD_1_PCOUT(27),
  PCOUT(28) => R1IN_4_4_ADD_1_PCOUT(28),
  PCOUT(29) => R1IN_4_4_ADD_1_PCOUT(29),
  PCOUT(30) => R1IN_4_4_ADD_1_PCOUT(30),
  PCOUT(31) => R1IN_4_4_ADD_1_PCOUT(31),
  PCOUT(32) => R1IN_4_4_ADD_1_PCOUT(32),
  PCOUT(33) => R1IN_4_4_ADD_1_PCOUT(33),
  PCOUT(34) => R1IN_4_4_ADD_1_PCOUT(34),
  PCOUT(35) => R1IN_4_4_ADD_1_PCOUT(35),
  PCOUT(36) => R1IN_4_4_ADD_1_PCOUT(36),
  PCOUT(37) => R1IN_4_4_ADD_1_PCOUT(37),
  PCOUT(38) => R1IN_4_4_ADD_1_PCOUT(38),
  PCOUT(39) => R1IN_4_4_ADD_1_PCOUT(39),
  PCOUT(40) => R1IN_4_4_ADD_1_PCOUT(40),
  PCOUT(41) => R1IN_4_4_ADD_1_PCOUT(41),
  PCOUT(42) => R1IN_4_4_ADD_1_PCOUT(42),
  PCOUT(43) => R1IN_4_4_ADD_1_PCOUT(43),
  PCOUT(44) => R1IN_4_4_ADD_1_PCOUT(44),
  PCOUT(45) => R1IN_4_4_ADD_1_PCOUT(45),
  PCOUT(46) => R1IN_4_4_ADD_1_PCOUT(46),
  PCOUT(47) => R1IN_4_4_ADD_1_PCOUT(47));
II_GND: GND port map (
    G => NN_1);
II_VCC: VCC port map (
    P => NN_2);
PRODUCT(17) <= NN_11;
end beh;

