-- Gaisler Ethernet core
  constant CFG_GRETH2 	 : integer := CONFIG_GRETH2_ENABLE;
  constant CFG_GRETH21G	 : integer := CONFIG_GRETH2_GIGA;
  constant CFG_ETH2_FIFO : integer := CFG_GRETH2_FIFO;

