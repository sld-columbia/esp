../ariane/ariane/src/register_interface/src/apb_to_reg.sv