../ariane/riscv_plic_apb_wrap.vhd