-- Second JTAG based DSU interface
  constant CFG_AHB_JTAG2	: integer := CONFIG_DSU_JTAG2;

