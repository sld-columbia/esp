library ieee;
use ieee.std_logic_1164.all;

package pads_loc is

  constant clk_div_acc0_pad_loc : std_logic := '0';
  constant clk_div_acc1_pad_loc : std_logic := '0';
  constant clk_div_cpu_pad_loc : std_logic := '0';
  constant dummy_pad_loc : std_logic := '0';
  constant erx_clk_pad_loc : std_logic := '0';
  constant erxd_pad_loc : std_logic_vector(3 downto 0) := "0000";
  constant erx_dv_pad_loc : std_logic := '0';
  constant etx_clk_pad_loc : std_logic := '0';
  constant ext_clk_acc0_pad_loc : std_logic := '0';
  constant ext_clk_acc1_pad_loc : std_logic := '0';
  constant ext_clk_cpu_pad_loc : std_logic := '0';
  constant fpga_clk_in_pad_loc : std_logic_vector(3 downto 0) := "0011";
  constant fpga_clk_out_pad_loc : std_logic_vector(3 downto 0) := "0011";
  constant fpga_credit_in_pad_loc : std_logic_vector(3 downto 0) := "0011";
  constant fpga_credit_out_pad_loc : std_logic_vector(3 downto 0) := "0011";
  constant fpga_data_pad_loc : std_logic_vector(255 downto 0) := "1111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000";
  constant fpga_valid_in_pad_loc : std_logic_vector(3 downto 0) := "0111";
  constant fpga_valid_out_pad_loc : std_logic_vector(3 downto 0) := "0111";
  constant lpddr0_addr_pad_loc : std_logic_vector(15 downto 0) := "0000000000000000";
  constant lpddr0_ba_pad_loc : std_logic_vector(2 downto 0) := "000";
  constant lpddr0_cas_n_pad_loc : std_logic := '0';
  constant lpddr0_cke_pad_loc : std_logic := '0';
  constant lpddr0_ck_n_pad_loc : std_logic := '0';
  constant lpddr0_ck_p_pad_loc : std_logic := '0';
  constant lpddr0_cs_n_pad_loc : std_logic := '0';
  constant lpddr0_dm_pad_loc : std_logic_vector(3 downto 0) := "0000";
  constant lpddr0_dq_pad_loc : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
  constant lpddr0_dqs_n_pad_loc : std_logic_vector(3 downto 0) := "0000";
  constant lpddr0_dqs_p_pad_loc : std_logic_vector(3 downto 0) := "0000";
  constant lpddr0_odt_pad_loc : std_logic := '0';
  constant lpddr0_ras_n_pad_loc : std_logic := '0';
  constant lpddr0_reset_n_pad_loc : std_logic := '0';
  constant lpddr0_we_n_pad_loc : std_logic := '0';
  constant reset_pad_loc : std_logic := '0';
  constant reset_o2_pad_loc : std_logic := '0';
  constant tclk_pad_loc : std_logic := '0';
  constant tdi_acc2_pad_loc : std_logic := '0';
  constant tdi_acc3_pad_loc : std_logic := '0';
  constant tdi_acc6_pad_loc : std_logic := '0';
  constant tdi_acc7_pad_loc : std_logic := '0';
  constant tdi_cpu_pad_loc : std_logic := '0';
  constant tdo_acc2_pad_loc : std_logic := '0';
  constant tdo_acc3_pad_loc : std_logic := '0';
  constant tdo_acc6_pad_loc : std_logic := '0';
  constant tdo_acc7_pad_loc : std_logic := '0';
  constant tdo_cpu_pad_loc : std_logic := '0';
  constant tms_pad_loc : std_logic := '0';
  constant unused_pad_loc : std_logic := '0';
  constant ivr_avs_clk_pad_loc : std_logic := '0';
  constant ivr_avs_dat_pad_loc : std_logic := '0';
  constant ivr_avs_sdat_pad_loc : std_logic := '0';
  constant ivr_control_pad_loc : std_logic := '0';
  constant clk_div_io_pad_loc : std_logic := '1';
  constant clk_div_mem_pad_loc : std_logic := '1';
  constant clk_div_noc_pad_loc : std_logic := '1';
  constant emdc_pad_loc : std_logic := '1';
  constant emdio_pad_loc : std_logic := '1';
  constant erx_col_pad_loc : std_logic := '1';
  constant erx_crs_pad_loc : std_logic := '1';
  constant erx_er_pad_loc : std_logic := '1';
  constant etxd_pad_loc : std_logic_vector(3 downto 0) := "1111";
  constant etx_en_pad_loc : std_logic := '1';
  constant etx_er_pad_loc : std_logic := '1';
  constant ext_clk_io_pad_loc : std_logic := '1';
  constant ext_clk_mem_pad_loc : std_logic := '1';
  constant ext_clk_noc_pad_loc : std_logic := '1';
  constant lpddr1_addr_pad_loc : std_logic_vector(15 downto 0) := "1111111111111111";
  constant lpddr1_ba_pad_loc : std_logic_vector(2 downto 0) := "111";
  constant lpddr1_cas_n_pad_loc : std_logic := '1';
  constant lpddr1_cke_pad_loc : std_logic := '1';
  constant lpddr1_ck_n_pad_loc : std_logic := '1';
  constant lpddr1_ck_p_pad_loc : std_logic := '1';
  constant lpddr1_cs_n_pad_loc : std_logic := '1';
  constant lpddr1_dm_pad_loc : std_logic_vector(3 downto 0) := "1111";
  constant lpddr1_dq_pad_loc : std_logic_vector(31 downto 0) := "11111111111111111111111111111111";
  constant lpddr1_dqs_n_pad_loc : std_logic_vector(3 downto 0) := "1111";
  constant lpddr1_dqs_p_pad_loc : std_logic_vector(3 downto 0) := "1111";
  constant lpddr1_odt_pad_loc : std_logic := '1';
  constant lpddr1_ras_n_pad_loc : std_logic := '1';
  constant lpddr1_reset_n_pad_loc : std_logic := '1';
  constant lpddr1_we_n_pad_loc : std_logic := '1';
  constant tdi_acc0_pad_loc : std_logic := '1';
  constant tdi_acc1_pad_loc : std_logic := '1';
  constant tdi_acc4_pad_loc : std_logic := '1';
  constant tdi_acc5_pad_loc : std_logic := '1';
  constant tdi_io_pad_loc : std_logic := '1';
  constant tdi_mem_pad_loc : std_logic := '1';
  constant tdo_acc0_pad_loc : std_logic := '1';
  constant tdo_acc1_pad_loc : std_logic := '1';
  constant tdo_acc4_pad_loc : std_logic := '1';
  constant tdo_acc5_pad_loc : std_logic := '1';
  constant tdo_io_pad_loc : std_logic := '1';
  constant tdo_mem_pad_loc : std_logic := '1';
  constant uart_ctsn_pad_loc : std_logic := '1';
  constant uart_rtsn_pad_loc : std_logic := '1';
  constant uart_rxd_pad_loc : std_logic := '1';
  constant uart_txd_pad_loc : std_logic := '1';
  constant ivr_gpio_pad_loc : std_logic_vector(3 downto 0) := "1111";
  constant ivr_pmb_dat_pad_loc : std_logic := '1';
  constant ivr_pmb_clk_pad_loc : std_logic := '1';

end package pads_loc;
