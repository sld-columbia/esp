-- AMBA System ACE Interface Controller
  constant CFG_GRACECTRL : integer := CONFIG_GRACECTRL;

