../vortex/hw/rtl/VX_scope.vh