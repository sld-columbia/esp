-- I2C to AHB bridge
  constant CFG_I2C2AHB         : integer := CONFIG_I2C2AHB;
  constant CFG_I2C2AHB_APB     : integer := CONFIG_I2C2AHB_APB;
  constant CFG_I2C2AHB_ADDRH   : integer := 16#CONFIG_I2C2AHB_ADDRH#;
  constant CFG_I2C2AHB_ADDRL   : integer := 16#CONFIG_I2C2AHB_ADDRL#;
  constant CFG_I2C2AHB_MASKH   : integer := 16#CONFIG_I2C2AHB_MASKH#;
  constant CFG_I2C2AHB_MASKL   : integer := 16#CONFIG_I2C2AHB_MASKL#;
  constant CFG_I2C2AHB_RESEN   : integer := CONFIG_I2C2AHB_RESEN;
  constant CFG_I2C2AHB_SADDR   : integer := 16#CONFIG_I2C2AHB_SADDR#;
  constant CFG_I2C2AHB_CADDR   : integer := 16#CONFIG_I2C2AHB_CADDR#;
  constant CFG_I2C2AHB_FILTER  : integer := CONFIG_I2C2AHB_FILTER;

