../vortex/hw/rtl/VX_platform.vh