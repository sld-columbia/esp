../vortex/hw/dpi/util_dpi.vh