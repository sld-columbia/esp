../vortex/hw/rtl/VX_config.vh