../../../../rtl/cores/ariane/ariane/src/fpu/src/fpnew_pkg.sv