../vortex/hw/rtl/fp_cores/VX_fpu_types.vh