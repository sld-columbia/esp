-- Second GPIO port
  constant CFG_GRGPIO2_ENABLE : integer := CONFIG_GRGPIO2_ENABLE;
  constant CFG_GRGPIO2_IMASK  : integer := 16#CONFIG_GRGPIO2_IMASK#;
  constant CFG_GRGPIO2_WIDTH  : integer := CONFIG_GRGPIO2_WIDTH;

