../ariane/ariane/src/register_interface/src/reg_intf.sv