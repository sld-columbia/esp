-- VGA and PS2/ interface
  constant CFG_KBD_ENABLE  : integer := CONFIG_KBD_ENABLE;
  constant CFG_VGA_ENABLE  : integer := CONFIG_VGA_ENABLE;
  constant CFG_SVGA_ENABLE : integer := CONFIG_SVGA_ENABLE;
  constant CFG_SVGA_MEMORY_HADDR : integer := 16#CONFIG_SVGA_MEMORY_HADDR#;

