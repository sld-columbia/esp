-- FT AHB RAM
  constant CFG_FTAHBRAM_EN       : integer := CONFIG_FTAHBRAM_ENABLE;
  constant CFG_FTAHBRAM_SZ       : integer := CONFIG_FTAHBRAM_SZ;
  constant CFG_FTAHBRAM_ADDR     : integer := 16#CONFIG_FTAHBRAM_START#;
  constant CFG_FTAHBRAM_PIPE     : integer := CONFIG_FTAHBRAM_PIPE;
  constant CFG_FTAHBRAM_EDAC     : integer := CONFIG_FTAHBRAM_EDAC;
  constant CFG_FTAHBRAM_SCRU     : integer := CONFIG_FTAHBRAM_AUTOSCRUB;
  constant CFG_FTAHBRAM_ECNT     : integer := CONFIG_FTAHBRAM_ERRORCNTR;
  constant CFG_FTAHBRAM_EBIT     : integer := CONFIG_FTAHBRAM_CNTBITS;

