rtl/fp_cores/xilinx/vc707/acl_fdiv/acl_fdiv.ip_user_files/ipstatic/hdl/axi_utils_v2_0_vh_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fdiv/acl_fdiv.ip_user_files/ipstatic/hdl/floating_point_v7_1_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fdiv/acl_fdiv.ip_user_files/ipstatic/hdl/mult_gen_v12_0_vh_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fdiv/acl_fdiv.ip_user_files/ipstatic/hdl/xbip_bram18k_v3_0_vh_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fdiv/acl_fdiv.ip_user_files/ipstatic/hdl/xbip_dsp48_addsub_v3_0_vh_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fdiv/acl_fdiv.ip_user_files/ipstatic/hdl/xbip_dsp48_multadd_v3_0_vh_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fdiv/acl_fdiv.ip_user_files/ipstatic/hdl/xbip_dsp48_wrapper_v3_0_vh_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fdiv/acl_fdiv.ip_user_files/ipstatic/hdl/xbip_pipe_v3_0_vh_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fdiv/acl_fdiv.ip_user_files/ipstatic/hdl/xbip_utils_v3_0_vh_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fsqrt/acl_fsqrt.ip_user_files/ipstatic/hdl/axi_utils_v2_0_vh_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fsqrt/acl_fsqrt.ip_user_files/ipstatic/hdl/floating_point_v7_1_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fsqrt/acl_fsqrt.ip_user_files/ipstatic/hdl/mult_gen_v12_0_vh_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fsqrt/acl_fsqrt.ip_user_files/ipstatic/hdl/xbip_bram18k_v3_0_vh_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fsqrt/acl_fsqrt.ip_user_files/ipstatic/hdl/xbip_dsp48_addsub_v3_0_vh_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fsqrt/acl_fsqrt.ip_user_files/ipstatic/hdl/xbip_dsp48_multadd_v3_0_vh_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fsqrt/acl_fsqrt.ip_user_files/ipstatic/hdl/xbip_dsp48_wrapper_v3_0_vh_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fsqrt/acl_fsqrt.ip_user_files/ipstatic/hdl/xbip_pipe_v3_0_vh_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fsqrt/acl_fsqrt.ip_user_files/ipstatic/hdl/xbip_utils_v3_0_vh_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fmadd/acl_fmadd.ip_user_files/ipstatic/hdl/axi_utils_v2_0_vh_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fmadd/acl_fmadd.ip_user_files/ipstatic/hdl/floating_point_v7_1_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fmadd/acl_fmadd.ip_user_files/ipstatic/hdl/mult_gen_v12_0_vh_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fmadd/acl_fmadd.ip_user_files/ipstatic/hdl/xbip_bram18k_v3_0_vh_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fmadd/acl_fmadd.ip_user_files/ipstatic/hdl/xbip_dsp48_addsub_v3_0_vh_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fmadd/acl_fmadd.ip_user_files/ipstatic/hdl/xbip_dsp48_multadd_v3_0_vh_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fmadd/acl_fmadd.ip_user_files/ipstatic/hdl/xbip_dsp48_wrapper_v3_0_vh_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fmadd/acl_fmadd.ip_user_files/ipstatic/hdl/xbip_pipe_v3_0_vh_rfs.vhd
rtl/fp_cores/xilinx/vc707/acl_fmadd/acl_fmadd.ip_user_files/ipstatic/hdl/xbip_utils_v3_0_vh_rfs.vhd
