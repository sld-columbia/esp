../vortex/hw/rtl/VX_trace_instr.vh