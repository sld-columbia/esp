-- Copyright (c) 2011-2024 Columbia University, System Level Design Group
-- SPDX-License-Identifier: Apache-2.0

-----------------------------------------------------------------------------
--  Accelerator Tile
------------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;
  use work.esp_global.all;
  use work.amba.all;
  use work.stdlib.all;
  use work.sld_devices.all;
  use work.devices.all;
  use work.gencomp.all;
  use work.monitor_pkg.all;
  use work.esp_csr_pkg.all;
  use work.jtag_pkg.all;
  use work.sldacc.all;
  use work.nocpackage.all;
  use work.cachepackage.all;
  use work.tile.all;
  use work.misc.all;
  use work.coretypes.all;
  use work.esp_acc_regmap.all;
  use work.socmap.all;
  use work.grlib_config.all;
  use work.tiles_pkg.all;

entity asic_tile_acc is
  generic (
    this_hls_conf : hlscfg_t             := 0;
    this_device   : devid_t              := 0;
    this_irq_type : integer              := 0;
    this_has_l2   : integer range 0 to 1 := 0;
    has_sync      : integer range 0 to 1 := 1;
    router_ports  : ports_vec            := "11111";
    this_has_dco  : integer range 0 to 1 := 0
  );
  port (
    rst          : in    std_ulogic;
    sys_clk      : in    std_ulogic; -- NoC clock
    sys_clk_lock : in    std_ulogic; -- sys_clk_lock
    ext_clk      : in    std_ulogic; -- backup tile clock
    clk_div      : out   std_ulogic; -- tile clock monitor for testing purposes
    -- Test interface
    tdi  : in    std_logic;
    tdo  : out   std_logic;
    tms  : in    std_logic;
    tclk : in    std_logic;
    -- Pad configuratio
    pad_cfg : out   std_logic_vector(ESP_CSR_PAD_CFG_MSB - ESP_CSR_PAD_CFG_LSB downto 0);
    -- NOC
    noc1_data_n_in     : in    coh_noc_flit_type;
    noc1_data_s_in     : in    coh_noc_flit_type;
    noc1_data_w_in     : in    coh_noc_flit_type;
    noc1_data_e_in     : in    coh_noc_flit_type;
    noc1_data_void_in  : in    std_logic_vector(3 downto 0);
    noc1_stop_in       : in    std_logic_vector(3 downto 0);
    noc1_data_n_out    : out   coh_noc_flit_type;
    noc1_data_s_out    : out   coh_noc_flit_type;
    noc1_data_w_out    : out   coh_noc_flit_type;
    noc1_data_e_out    : out   coh_noc_flit_type;
    noc1_data_void_out : out   std_logic_vector(3 downto 0);
    noc1_stop_out      : out   std_logic_vector(3 downto 0);
    noc2_data_n_in     : in    coh_noc_flit_type;
    noc2_data_s_in     : in    coh_noc_flit_type;
    noc2_data_w_in     : in    coh_noc_flit_type;
    noc2_data_e_in     : in    coh_noc_flit_type;
    noc2_data_void_in  : in    std_logic_vector(3 downto 0);
    noc2_stop_in       : in    std_logic_vector(3 downto 0);
    noc2_data_n_out    : out   coh_noc_flit_type;
    noc2_data_s_out    : out   coh_noc_flit_type;
    noc2_data_w_out    : out   coh_noc_flit_type;
    noc2_data_e_out    : out   coh_noc_flit_type;
    noc2_data_void_out : out   std_logic_vector(3 downto 0);
    noc2_stop_out      : out   std_logic_vector(3 downto 0);
    noc3_data_n_in     : in    coh_noc_flit_type;
    noc3_data_s_in     : in    coh_noc_flit_type;
    noc3_data_w_in     : in    coh_noc_flit_type;
    noc3_data_e_in     : in    coh_noc_flit_type;
    noc3_data_void_in  : in    std_logic_vector(3 downto 0);
    noc3_stop_in       : in    std_logic_vector(3 downto 0);
    noc3_data_n_out    : out   coh_noc_flit_type;
    noc3_data_s_out    : out   coh_noc_flit_type;
    noc3_data_w_out    : out   coh_noc_flit_type;
    noc3_data_e_out    : out   coh_noc_flit_type;
    noc3_data_void_out : out   std_logic_vector(3 downto 0);
    noc3_stop_out      : out   std_logic_vector(3 downto 0);
    noc4_data_n_in     : in    dma_noc_flit_type;
    noc4_data_s_in     : in    dma_noc_flit_type;
    noc4_data_w_in     : in    dma_noc_flit_type;
    noc4_data_e_in     : in    dma_noc_flit_type;
    noc4_data_void_in  : in    std_logic_vector(3 downto 0);
    noc4_stop_in       : in    std_logic_vector(3 downto 0);
    noc4_data_n_out    : out   dma_noc_flit_type;
    noc4_data_s_out    : out   dma_noc_flit_type;
    noc4_data_w_out    : out   dma_noc_flit_type;
    noc4_data_e_out    : out   dma_noc_flit_type;
    noc4_data_void_out : out   std_logic_vector(3 downto 0);
    noc4_stop_out      : out   std_logic_vector(3 downto 0);
    noc5_data_n_in     : in    misc_noc_flit_type;
    noc5_data_s_in     : in    misc_noc_flit_type;
    noc5_data_w_in     : in    misc_noc_flit_type;
    noc5_data_e_in     : in    misc_noc_flit_type;
    noc5_data_void_in  : in    std_logic_vector(3 downto 0);
    noc5_stop_in       : in    std_logic_vector(3 downto 0);
    noc5_data_n_out    : out   misc_noc_flit_type;
    noc5_data_s_out    : out   misc_noc_flit_type;
    noc5_data_w_out    : out   misc_noc_flit_type;
    noc5_data_e_out    : out   misc_noc_flit_type;
    noc5_data_void_out : out   std_logic_vector(3 downto 0);
    noc5_stop_out      : out   std_logic_vector(3 downto 0);
    noc6_data_n_in     : in    dma_noc_flit_type;
    noc6_data_s_in     : in    dma_noc_flit_type;
    noc6_data_w_in     : in    dma_noc_flit_type;
    noc6_data_e_in     : in    dma_noc_flit_type;
    noc6_data_void_in  : in    std_logic_vector(3 downto 0);
    noc6_stop_in       : in    std_logic_vector(3 downto 0);
    noc6_data_n_out    : out   dma_noc_flit_type;
    noc6_data_s_out    : out   dma_noc_flit_type;
    noc6_data_w_out    : out   dma_noc_flit_type;
    noc6_data_e_out    : out   dma_noc_flit_type;
    noc6_data_void_out : out   std_logic_vector(3 downto 0);
    noc6_stop_out      : out   std_logic_vector(3 downto 0)
  );
end entity asic_tile_acc;

architecture rtl of asic_tile_acc is

  constant EXT_CLK_SEL_DEFAULT : std_ulogic := '0';

  -- Tile clock and reset (only for I/O tile)
  signal raw_rstn : std_ulogic;
  signal dco_clk  : std_ulogic;
  signal dco_rstn : std_ulogic;
  signal tile_rst : std_ulogic;
  --  signal dco_clk_lock : std_ulogic;

  -- Tile parameters
  signal this_local_y : local_yx;
  signal this_local_x : local_yx;

  -- Tile interface signals
  signal test_rstn             : std_ulogic;
  signal test1_output_port_s   : coh_noc_flit_type;
  signal test1_data_void_out_s : std_ulogic;
  signal test1_stop_in_s       : std_ulogic;
  signal test2_output_port_s   : coh_noc_flit_type;
  signal test2_data_void_out_s : std_ulogic;
  signal test2_stop_in_s       : std_ulogic;
  signal test3_output_port_s   : coh_noc_flit_type;
  signal test3_data_void_out_s : std_ulogic;
  signal test3_stop_in_s       : std_ulogic;
  signal test4_output_port_s   : dma_noc_flit_type;
  signal test4_data_void_out_s : std_ulogic;
  signal test4_stop_in_s       : std_ulogic;
  signal test5_output_port_s   : misc_noc_flit_type;
  signal test5_data_void_out_s : std_ulogic;
  signal test5_stop_in_s       : std_ulogic;
  signal test6_output_port_s   : dma_noc_flit_type;
  signal test6_data_void_out_s : std_ulogic;
  signal test6_stop_in_s       : std_ulogic;
  signal test1_input_port_s    : coh_noc_flit_type;
  signal test1_data_void_in_s  : std_ulogic;
  signal test1_stop_out_s      : std_ulogic;
  signal test2_input_port_s    : coh_noc_flit_type;
  signal test2_data_void_in_s  : std_ulogic;
  signal test2_stop_out_s      : std_ulogic;
  signal test3_input_port_s    : coh_noc_flit_type;
  signal test3_data_void_in_s  : std_ulogic;
  signal test3_stop_out_s      : std_ulogic;
  signal test4_input_port_s    : dma_noc_flit_type;
  signal test4_data_void_in_s  : std_ulogic;
  signal test4_stop_out_s      : std_ulogic;
  signal test5_input_port_s    : misc_noc_flit_type;
  signal test5_data_void_in_s  : std_ulogic;
  signal test5_stop_out_s      : std_ulogic;
  signal test6_input_port_s    : dma_noc_flit_type;
  signal test6_data_void_in_s  : std_ulogic;
  signal test6_stop_out_s      : std_ulogic;

  signal noc1_mon_noc_vec_int : monitor_noc_type;
  signal noc2_mon_noc_vec_int : monitor_noc_type;
  signal noc3_mon_noc_vec_int : monitor_noc_type;
  signal noc4_mon_noc_vec_int : monitor_noc_type;
  signal noc5_mon_noc_vec_int : monitor_noc_type;
  signal noc6_mon_noc_vec_int : monitor_noc_type;

  -- Noc signals
  signal noc_rstn               : std_ulogic;
  signal noc1_stop_in_s         : std_logic_vector(4 downto 0);
  signal noc1_stop_out_s        : std_logic_vector(4 downto 0);
  signal noc1_acc_stop_in       : std_ulogic;
  signal noc1_acc_stop_out      : std_ulogic;
  signal noc1_data_void_in_s    : std_logic_vector(4 downto 0);
  signal noc1_data_void_out_s   : std_logic_vector(4 downto 0);
  signal noc1_acc_data_void_in  : std_ulogic;
  signal noc1_acc_data_void_out : std_ulogic;
  signal noc2_stop_in_s         : std_logic_vector(4 downto 0);
  signal noc2_stop_out_s        : std_logic_vector(4 downto 0);
  signal noc2_acc_stop_in       : std_ulogic;
  signal noc2_acc_stop_out      : std_ulogic;
  signal noc2_data_void_in_s    : std_logic_vector(4 downto 0);
  signal noc2_data_void_out_s   : std_logic_vector(4 downto 0);
  signal noc2_acc_data_void_in  : std_ulogic;
  signal noc2_acc_data_void_out : std_ulogic;
  signal noc3_stop_in_s         : std_logic_vector(4 downto 0);
  signal noc3_stop_out_s        : std_logic_vector(4 downto 0);
  signal noc3_acc_stop_in       : std_ulogic;
  signal noc3_acc_stop_out      : std_ulogic;
  signal noc3_data_void_in_s    : std_logic_vector(4 downto 0);
  signal noc3_data_void_out_s   : std_logic_vector(4 downto 0);
  signal noc3_acc_data_void_in  : std_ulogic;
  signal noc3_acc_data_void_out : std_ulogic;
  signal noc4_stop_in_s         : std_logic_vector(4 downto 0);
  signal noc4_stop_out_s        : std_logic_vector(4 downto 0);
  signal noc4_acc_stop_in       : std_ulogic;
  signal noc4_acc_stop_out      : std_ulogic;
  signal noc4_data_void_in_s    : std_logic_vector(4 downto 0);
  signal noc4_data_void_out_s   : std_logic_vector(4 downto 0);
  signal noc4_acc_data_void_in  : std_ulogic;
  signal noc4_acc_data_void_out : std_ulogic;
  signal noc5_stop_in_s         : std_logic_vector(4 downto 0);
  signal noc5_stop_out_s        : std_logic_vector(4 downto 0);
  signal noc5_acc_stop_in       : std_ulogic;
  signal noc5_acc_stop_out      : std_ulogic;
  signal noc5_data_void_in_s    : std_logic_vector(4 downto 0);
  signal noc5_data_void_out_s   : std_logic_vector(4 downto 0);
  signal noc5_acc_data_void_in  : std_ulogic;
  signal noc5_acc_data_void_out : std_ulogic;
  signal noc6_stop_in_s         : std_logic_vector(4 downto 0);
  signal noc6_stop_out_s        : std_logic_vector(4 downto 0);
  signal noc6_acc_stop_in       : std_ulogic;
  signal noc6_acc_stop_out      : std_ulogic;
  signal noc6_data_void_in_s    : std_logic_vector(4 downto 0);
  signal noc6_data_void_out_s   : std_logic_vector(4 downto 0);
  signal noc6_acc_data_void_in  : std_ulogic;
  signal noc6_acc_data_void_out : std_ulogic;
  signal noc1_input_port        : coh_noc_flit_type;
  signal noc2_input_port        : coh_noc_flit_type;
  signal noc3_input_port        : coh_noc_flit_type;
  signal noc4_input_port        : dma_noc_flit_type;
  signal noc5_input_port        : misc_noc_flit_type;
  signal noc6_input_port        : dma_noc_flit_type;
  signal noc1_output_port       : coh_noc_flit_type;
  signal noc2_output_port       : coh_noc_flit_type;
  signal noc3_output_port       : coh_noc_flit_type;
  signal noc4_output_port       : dma_noc_flit_type;
  signal noc5_output_port       : misc_noc_flit_type;
  signal noc6_output_port       : dma_noc_flit_type;

  attribute keep              : string;
  attribute keep of noc1_acc_stop_in       : signal is "true";
  attribute keep of noc1_acc_stop_out      : signal is "true";
  attribute keep of noc1_acc_data_void_in  : signal is "true";
  attribute keep of noc1_acc_data_void_out : signal is "true";
  attribute keep of noc1_input_port        : signal is "true";
  attribute keep of noc1_output_port       : signal is "true";
  attribute keep of noc1_data_n_in         : signal is "true";
  attribute keep of noc1_data_s_in         : signal is "true";
  attribute keep of noc1_data_w_in         : signal is "true";
  attribute keep of noc1_data_e_in         : signal is "true";
  attribute keep of noc1_data_void_in      : signal is "true";
  attribute keep of noc1_stop_in           : signal is "true";
  attribute keep of noc1_data_n_out        : signal is "true";
  attribute keep of noc1_data_s_out        : signal is "true";
  attribute keep of noc1_data_w_out        : signal is "true";
  attribute keep of noc1_data_e_out        : signal is "true";
  attribute keep of noc1_data_void_out     : signal is "true";
  attribute keep of noc1_stop_out          : signal is "true";
  attribute keep of noc2_acc_stop_in       : signal is "true";
  attribute keep of noc2_acc_stop_out      : signal is "true";
  attribute keep of noc2_acc_data_void_in  : signal is "true";
  attribute keep of noc2_acc_data_void_out : signal is "true";
  attribute keep of noc2_input_port        : signal is "true";
  attribute keep of noc2_output_port       : signal is "true";
  attribute keep of noc2_data_n_in         : signal is "true";
  attribute keep of noc2_data_s_in         : signal is "true";
  attribute keep of noc2_data_w_in         : signal is "true";
  attribute keep of noc2_data_e_in         : signal is "true";
  attribute keep of noc2_data_void_in      : signal is "true";
  attribute keep of noc2_stop_in           : signal is "true";
  attribute keep of noc2_data_n_out        : signal is "true";
  attribute keep of noc2_data_s_out        : signal is "true";
  attribute keep of noc2_data_w_out        : signal is "true";
  attribute keep of noc2_data_e_out        : signal is "true";
  attribute keep of noc2_data_void_out     : signal is "true";
  attribute keep of noc2_stop_out          : signal is "true";
  attribute keep of noc3_acc_stop_in       : signal is "true";
  attribute keep of noc3_acc_stop_out      : signal is "true";
  attribute keep of noc3_acc_data_void_in  : signal is "true";
  attribute keep of noc3_acc_data_void_out : signal is "true";
  attribute keep of noc3_input_port        : signal is "true";
  attribute keep of noc3_output_port       : signal is "true";
  attribute keep of noc3_data_n_in         : signal is "true";
  attribute keep of noc3_data_s_in         : signal is "true";
  attribute keep of noc3_data_w_in         : signal is "true";
  attribute keep of noc3_data_e_in         : signal is "true";
  attribute keep of noc3_data_void_in      : signal is "true";
  attribute keep of noc3_stop_in           : signal is "true";
  attribute keep of noc3_data_n_out        : signal is "true";
  attribute keep of noc3_data_s_out        : signal is "true";
  attribute keep of noc3_data_w_out        : signal is "true";
  attribute keep of noc3_data_e_out        : signal is "true";
  attribute keep of noc3_data_void_out     : signal is "true";
  attribute keep of noc3_stop_out          : signal is "true";
  attribute keep of noc4_acc_stop_in       : signal is "true";
  attribute keep of noc4_acc_stop_out      : signal is "true";
  attribute keep of noc4_acc_data_void_in  : signal is "true";
  attribute keep of noc4_acc_data_void_out : signal is "true";
  attribute keep of noc4_input_port        : signal is "true";
  attribute keep of noc4_output_port       : signal is "true";
  attribute keep of noc4_data_n_in         : signal is "true";
  attribute keep of noc4_data_s_in         : signal is "true";
  attribute keep of noc4_data_w_in         : signal is "true";
  attribute keep of noc4_data_e_in         : signal is "true";
  attribute keep of noc4_data_void_in      : signal is "true";
  attribute keep of noc4_stop_in           : signal is "true";
  attribute keep of noc4_data_n_out        : signal is "true";
  attribute keep of noc4_data_s_out        : signal is "true";
  attribute keep of noc4_data_w_out        : signal is "true";
  attribute keep of noc4_data_e_out        : signal is "true";
  attribute keep of noc4_data_void_out     : signal is "true";
  attribute keep of noc4_stop_out          : signal is "true";
  attribute keep of noc5_acc_stop_in       : signal is "true";
  attribute keep of noc5_acc_stop_out      : signal is "true";
  attribute keep of noc5_acc_data_void_in  : signal is "true";
  attribute keep of noc5_acc_data_void_out : signal is "true";
  attribute keep of noc5_input_port        : signal is "true";
  attribute keep of noc5_output_port       : signal is "true";
  attribute keep of noc5_data_n_in         : signal is "true";
  attribute keep of noc5_data_s_in         : signal is "true";
  attribute keep of noc5_data_w_in         : signal is "true";
  attribute keep of noc5_data_e_in         : signal is "true";
  attribute keep of noc5_data_void_in      : signal is "true";
  attribute keep of noc5_stop_in           : signal is "true";
  attribute keep of noc5_data_n_out        : signal is "true";
  attribute keep of noc5_data_s_out        : signal is "true";
  attribute keep of noc5_data_w_out        : signal is "true";
  attribute keep of noc5_data_e_out        : signal is "true";
  attribute keep of noc5_data_void_out     : signal is "true";
  attribute keep of noc5_stop_out          : signal is "true";
  attribute keep of noc6_acc_stop_in       : signal is "true";
  attribute keep of noc6_acc_stop_out      : signal is "true";
  attribute keep of noc6_acc_data_void_in  : signal is "true";
  attribute keep of noc6_acc_data_void_out : signal is "true";
  attribute keep of noc6_input_port        : signal is "true";
  attribute keep of noc6_output_port       : signal is "true";
  attribute keep of noc6_data_n_in         : signal is "true";
  attribute keep of noc6_data_s_in         : signal is "true";
  attribute keep of noc6_data_w_in         : signal is "true";
  attribute keep of noc6_data_e_in         : signal is "true";
  attribute keep of noc6_data_void_in      : signal is "true";
  attribute keep of noc6_stop_in           : signal is "true";
  attribute keep of noc6_data_n_out        : signal is "true";
  attribute keep of noc6_data_s_out        : signal is "true";
  attribute keep of noc6_data_w_out        : signal is "true";
  attribute keep of noc6_data_e_out        : signal is "true";
  attribute keep of noc6_data_void_out     : signal is "true";
  attribute keep of noc6_stop_out          : signal is "true";

begin

  rst_noc : component rstgen
    generic map (
      acthigh => 1, syncin => 0
    )
    port map (
rst,
 sys_clk,
 sys_clk_lock,
 noc_rstn,
 raw_rstn
    );

  rst_jtag : component rstgen
    generic map (
      acthigh => 1, syncin => 0
    )
    port map (
rst,
 tclk,
 '1',
 test_rstn,
 open
    );

  has_dco_rst : if this_has_dco = 1 generate
    tile_rst <= rst;
  end generate has_dco_rst;

  no_dco_rst : if this_has_dco /= 1 generate
    tile_rst <= noc_rstn;
  end generate no_dco_rst;

  -----------------------------------------------------------------------------
  -- JTAG for single tile testing / bypass when test_if_en = 0
  -----------------------------------------------------------------------------
  jtag_test_i : component jtag_test
    generic map (
      test_if_en => CFG_JTAG_EN
    )
    port map (
      rst                 => test_rstn,
      refclk              => dco_clk,
      tile_rst            => dco_rstn,
      tdi                 => tdi,
      tdo                 => tdo,
      tms                 => tms,
      tclk                => tclk,
      noc1_output_port    => noc1_output_port,
      noc1_data_void_out  => noc1_acc_data_void_out,
      noc1_stop_in        => noc1_acc_stop_in,
      noc2_output_port    => noc2_output_port,
      noc2_data_void_out  => noc2_acc_data_void_out,
      noc2_stop_in        => noc2_acc_stop_in,
      noc3_output_port    => noc3_output_port,
      noc3_data_void_out  => noc3_acc_data_void_out,
      noc3_stop_in        => noc3_acc_stop_in,
      noc4_output_port    => noc4_output_port,
      noc4_data_void_out  => noc4_acc_data_void_out,
      noc4_stop_in        => noc4_acc_stop_in,
      noc5_output_port    => noc5_output_port,
      noc5_data_void_out  => noc5_acc_data_void_out,
      noc5_stop_in        => noc5_acc_stop_in,
      noc6_output_port    => noc6_output_port,
      noc6_data_void_out  => noc6_acc_data_void_out,
      noc6_stop_in        => noc6_acc_stop_in,
      test1_output_port   => test1_output_port_s,
      test1_data_void_out => test1_data_void_out_s,
      test1_stop_in       => test1_stop_in_s,
      test2_output_port   => test2_output_port_s,
      test2_data_void_out => test2_data_void_out_s,
      test2_stop_in       => test2_stop_in_s,
      test3_output_port   => test3_output_port_s,
      test3_data_void_out => test3_data_void_out_s,
      test3_stop_in       => test3_stop_in_s,
      test4_output_port   => test4_output_port_s,
      test4_data_void_out => test4_data_void_out_s,
      test4_stop_in       => test4_stop_in_s,
      test5_output_port   => test5_output_port_s,
      test5_data_void_out => test5_data_void_out_s,
      test5_stop_in       => test5_stop_in_s,
      test6_output_port   => test6_output_port_s,
      test6_data_void_out => test6_data_void_out_s,
      test6_stop_in       => test6_stop_in_s,
      test1_input_port    => test1_input_port_s,
      test1_data_void_in  => test1_data_void_in_s,
      test1_stop_out      => test1_stop_out_s,
      test2_input_port    => test2_input_port_s,
      test2_data_void_in  => test2_data_void_in_s,
      test2_stop_out      => test2_stop_out_s,
      test3_input_port    => test3_input_port_s,
      test3_data_void_in  => test3_data_void_in_s,
      test3_stop_out      => test3_stop_out_s,
      test4_input_port    => test4_input_port_s,
      test4_data_void_in  => test4_data_void_in_s,
      test4_stop_out      => test4_stop_out_s,
      test5_input_port    => test5_input_port_s,
      test5_data_void_in  => test5_data_void_in_s,
      test5_stop_out      => test5_stop_out_s,
      test6_input_port    => test6_input_port_s,
      test6_data_void_in  => test6_data_void_in_s,
      test6_stop_out      => test6_stop_out_s,
      noc1_input_port     => noc1_input_port,
      noc1_data_void_in   => noc1_acc_data_void_in,
      noc1_stop_out       => noc1_acc_stop_out,
      noc2_input_port     => noc2_input_port,
      noc2_data_void_in   => noc2_acc_data_void_in,
      noc2_stop_out       => noc2_acc_stop_out,
      noc3_input_port     => noc3_input_port,
      noc3_data_void_in   => noc3_acc_data_void_in,
      noc3_stop_out       => noc3_acc_stop_out,
      noc4_input_port     => noc4_input_port,
      noc4_data_void_in   => noc4_acc_data_void_in,
      noc4_stop_out       => noc4_acc_stop_out,
      noc5_input_port     => noc5_input_port,
      noc5_data_void_in   => noc5_acc_data_void_in,
      noc5_stop_out       => noc5_acc_stop_out,
      noc6_input_port     => noc6_input_port,
      noc6_data_void_in   => noc6_acc_data_void_in,
      noc6_stop_out       => noc6_acc_stop_out
    );

  -----------------------------------------------------------------------------
  -- NOC Connections
  ----------------------------------------------------------------------------
  noc1_stop_in_s         <= noc1_acc_stop_in & noc1_stop_in;
  noc1_stop_out          <= noc1_stop_out_s(3 downto 0);
  noc1_acc_stop_out      <= noc1_stop_out_s(4);
  noc1_data_void_in_s    <= noc1_acc_data_void_in & noc1_data_void_in;
  noc1_data_void_out     <= noc1_data_void_out_s(3 downto 0);
  noc1_acc_data_void_out <= noc1_data_void_out_s(4);
  noc2_stop_in_s         <= noc2_acc_stop_in & noc2_stop_in;
  noc2_stop_out          <= noc2_stop_out_s(3 downto 0);
  noc2_acc_stop_out      <= noc2_stop_out_s(4);
  noc2_data_void_in_s    <= noc2_acc_data_void_in & noc2_data_void_in;
  noc2_data_void_out     <= noc2_data_void_out_s(3 downto 0);
  noc2_acc_data_void_out <= noc2_data_void_out_s(4);
  noc3_stop_in_s         <= noc3_acc_stop_in & noc3_stop_in;
  noc3_stop_out          <= noc3_stop_out_s(3 downto 0);
  noc3_acc_stop_out      <= noc3_stop_out_s(4);
  noc3_data_void_in_s    <= noc3_acc_data_void_in & noc3_data_void_in;
  noc3_data_void_out     <= noc3_data_void_out_s(3 downto 0);
  noc3_acc_data_void_out <= noc3_data_void_out_s(4);
  noc4_stop_in_s         <= noc4_acc_stop_in & noc4_stop_in;
  noc4_stop_out          <= noc4_stop_out_s(3 downto 0);
  noc4_acc_stop_out      <= noc4_stop_out_s(4);
  noc4_data_void_in_s    <= noc4_acc_data_void_in & noc4_data_void_in;
  noc4_data_void_out     <= noc4_data_void_out_s(3 downto 0);
  noc4_acc_data_void_out <= noc4_data_void_out_s(4);
  noc5_stop_in_s         <= noc5_acc_stop_in & noc5_stop_in;
  noc5_stop_out          <= noc5_stop_out_s(3 downto 0);
  noc5_acc_stop_out      <= noc5_stop_out_s(4);
  noc5_data_void_in_s    <= noc5_acc_data_void_in & noc5_data_void_in;
  noc5_data_void_out     <= noc5_data_void_out_s(3 downto 0);
  noc5_acc_data_void_out <= noc5_data_void_out_s(4);
  noc6_stop_in_s         <= noc6_acc_stop_in & noc6_stop_in;
  noc6_stop_out          <= noc6_stop_out_s(3 downto 0);
  noc6_acc_stop_out      <= noc6_stop_out_s(4);
  noc6_data_void_in_s    <= noc6_acc_data_void_in & noc6_data_void_in;
  noc6_data_void_out     <= noc6_data_void_out_s(3 downto 0);
  noc6_acc_data_void_out <= noc6_data_void_out_s(4);

  sync_noc_set_acc : component sync_noc_set
    generic map (
      ports    => ROUTER_PORTS,
      has_sync => HAS_SYNC
    )
    port map (
      clk                => sys_clk,
      clk_tile           => dco_clk,
      rst                => noc_rstn,
      rst_tile           => dco_rstn,
      const_local_x      => this_local_x,
      const_local_y      => this_local_y,
      noc1_data_n_in     => noc1_data_n_in,
      noc1_data_s_in     => noc1_data_s_in,
      noc1_data_w_in     => noc1_data_w_in,
      noc1_data_e_in     => noc1_data_e_in,
      noc1_input_port    => noc1_input_port,
      noc1_data_void_in  => noc1_data_void_in_s,
      noc1_stop_in       => noc1_stop_in_s,
      noc1_data_n_out    => noc1_data_n_out,
      noc1_data_s_out    => noc1_data_s_out,
      noc1_data_w_out    => noc1_data_w_out,
      noc1_data_e_out    => noc1_data_e_out,
      noc1_output_port   => noc1_output_port,
      noc1_data_void_out => noc1_data_void_out_s,
      noc1_stop_out      => noc1_stop_out_s,
      noc2_data_n_in     => noc2_data_n_in,
      noc2_data_s_in     => noc2_data_s_in,
      noc2_data_w_in     => noc2_data_w_in,
      noc2_data_e_in     => noc2_data_e_in,
      noc2_input_port    => noc2_input_port,
      noc2_data_void_in  => noc2_data_void_in_s,
      noc2_stop_in       => noc2_stop_in_s,
      noc2_data_n_out    => noc2_data_n_out,
      noc2_data_s_out    => noc2_data_s_out,
      noc2_data_w_out    => noc2_data_w_out,
      noc2_data_e_out    => noc2_data_e_out,
      noc2_output_port   => noc2_output_port,
      noc2_data_void_out => noc2_data_void_out_s,
      noc2_stop_out      => noc2_stop_out_s,
      noc3_data_n_in     => noc3_data_n_in,
      noc3_data_s_in     => noc3_data_s_in,
      noc3_data_w_in     => noc3_data_w_in,
      noc3_data_e_in     => noc3_data_e_in,
      noc3_input_port    => noc3_input_port,
      noc3_data_void_in  => noc3_data_void_in_s,
      noc3_stop_in       => noc3_stop_in_s,
      noc3_data_n_out    => noc3_data_n_out,
      noc3_data_s_out    => noc3_data_s_out,
      noc3_data_w_out    => noc3_data_w_out,
      noc3_data_e_out    => noc3_data_e_out,
      noc3_output_port   => noc3_output_port,
      noc3_data_void_out => noc3_data_void_out_s,
      noc3_stop_out      => noc3_stop_out_s,
      noc4_data_n_in     => noc4_data_n_in,
      noc4_data_s_in     => noc4_data_s_in,
      noc4_data_w_in     => noc4_data_w_in,
      noc4_data_e_in     => noc4_data_e_in,
      noc4_input_port    => noc4_input_port,
      noc4_data_void_in  => noc4_data_void_in_s,
      noc4_stop_in       => noc4_stop_in_s,
      noc4_data_n_out    => noc4_data_n_out,
      noc4_data_s_out    => noc4_data_s_out,
      noc4_data_w_out    => noc4_data_w_out,
      noc4_data_e_out    => noc4_data_e_out,
      noc4_output_port   => noc4_output_port,
      noc4_data_void_out => noc4_data_void_out_s,
      noc4_stop_out      => noc4_stop_out_s,
      noc5_data_n_in     => noc5_data_n_in,
      noc5_data_s_in     => noc5_data_s_in,
      noc5_data_w_in     => noc5_data_w_in,
      noc5_data_e_in     => noc5_data_e_in,
      noc5_input_port    => noc5_input_port,
      noc5_data_void_in  => noc5_data_void_in_s,
      noc5_stop_in       => noc5_stop_in_s,
      noc5_data_n_out    => noc5_data_n_out,
      noc5_data_s_out    => noc5_data_s_out,
      noc5_data_w_out    => noc5_data_w_out,
      noc5_data_e_out    => noc5_data_e_out,
      noc5_output_port   => noc5_output_port,
      noc5_data_void_out => noc5_data_void_out_s,
      noc5_stop_out      => noc5_stop_out_s,
      noc6_data_n_in     => noc6_data_n_in,
      noc6_data_s_in     => noc6_data_s_in,
      noc6_data_w_in     => noc6_data_w_in,
      noc6_data_e_in     => noc6_data_e_in,
      noc6_input_port    => noc6_input_port,
      noc6_data_void_in  => noc6_data_void_in_s,
      noc6_stop_in       => noc6_stop_in_s,
      noc6_data_n_out    => noc6_data_n_out,
      noc6_data_s_out    => noc6_data_s_out,
      noc6_data_w_out    => noc6_data_w_out,
      noc6_data_e_out    => noc6_data_e_out,
      noc6_output_port   => noc6_output_port,
      noc6_data_void_out => noc6_data_void_out_s,
      noc6_stop_out      => noc6_stop_out_s,
      noc1_mon_noc_vec   => noc1_mon_noc_vec_int,
      noc2_mon_noc_vec   => noc2_mon_noc_vec_int,
      noc3_mon_noc_vec   => noc3_mon_noc_vec_int,
      noc4_mon_noc_vec   => noc4_mon_noc_vec_int,
      noc5_mon_noc_vec   => noc5_mon_noc_vec_int,
      noc6_mon_noc_vec   => noc6_mon_noc_vec_int
    );

  tile_acc_1 : component tile_acc
    generic map (
      this_hls_conf      => this_hls_conf,
      this_device        => this_device,
      this_irq_type      => this_irq_type,
      this_has_l2        => this_has_l2,
      this_has_dvfs      => 0,
      this_has_pll       => 0,
      this_has_dco       => this_has_dco,
      this_extra_clk_buf => 0
    )
    port map (
      raw_rstn            => raw_rstn,
      tile_rst            => tile_rst,
      refclk              => ext_clk,
      pllbypass           => ext_clk_sel_default,
      pllclk              => clk_div,
      dco_clk             => dco_clk,
      dco_rstn            => dco_rstn,
      pad_cfg             => pad_cfg,
      local_x             => this_local_x,
      local_y             => this_local_y,
      test1_output_port   => test1_output_port_s,
      test1_data_void_out => test1_data_void_out_s,
      test1_stop_in       => test1_stop_out_s,
      test1_input_port    => test1_input_port_s,
      test1_data_void_in  => test1_data_void_in_s,
      test1_stop_out      => test1_stop_in_s,
      test2_output_port   => test2_output_port_s,
      test2_data_void_out => test2_data_void_out_s,
      test2_stop_in       => test2_stop_out_s,
      test2_input_port    => test2_input_port_s,
      test2_data_void_in  => test2_data_void_in_s,
      test2_stop_out      => test2_stop_in_s,
      test3_output_port   => test3_output_port_s,
      test3_data_void_out => test3_data_void_out_s,
      test3_stop_in       => test3_stop_out_s,
      test3_input_port    => test3_input_port_s,
      test3_data_void_in  => test3_data_void_in_s,
      test3_stop_out      => test3_stop_in_s,
      test4_output_port   => test4_output_port_s,
      test4_data_void_out => test4_data_void_out_s,
      test4_stop_in       => test4_stop_out_s,
      test4_input_port    => test4_input_port_s,
      test4_data_void_in  => test4_data_void_in_s,
      test4_stop_out      => test4_stop_in_s,
      test5_output_port   => test5_output_port_s,
      test5_data_void_out => test5_data_void_out_s,
      test5_stop_in       => test5_stop_out_s,
      test5_input_port    => test5_input_port_s,
      test5_data_void_in  => test5_data_void_in_s,
      test5_stop_out      => test5_stop_in_s,
      test6_output_port   => test6_output_port_s,
      test6_data_void_out => test6_data_void_out_s,
      test6_stop_in       => test6_stop_out_s,
      test6_input_port    => test6_input_port_s,
      test6_data_void_in  => test6_data_void_in_s,
      test6_stop_out      => test6_stop_in_s,
      noc1_mon_noc_vec    => noc1_mon_noc_vec_int,
      noc2_mon_noc_vec    => noc2_mon_noc_vec_int,
      noc3_mon_noc_vec    => noc3_mon_noc_vec_int,
      noc4_mon_noc_vec    => noc4_mon_noc_vec_int,
      noc5_mon_noc_vec    => noc5_mon_noc_vec_int,
      noc6_mon_noc_vec    => noc6_mon_noc_vec_int,
      mon_dvfs_in         => monitor_dvfs_none,
      mon_acc             => open,
      mon_cache           => open,
      mon_dvfs            => open
    );

end architecture rtl;
