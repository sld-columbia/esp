-- I2C slave
  constant CFG_I2CSLV_ENABLE   : integer := CONFIG_I2CSLV_ENABLE;
  constant CFG_I2CSLV_HARDADDR : integer := CONFIG_I2CSLV_HARDADDR;
  constant CFG_I2CSLV_TENBIT   : integer := CONFIG_I2CSLV_TENBIT;
  constant CFG_I2CSLV_I2CADDR  : integer := CONFIG_I2CSLV_I2CADDR;
  

