-- JTAG boundary-scan chain
  constant CFG_BOUNDSCAN_EN	: integer := CONFIG_BOUNDSCAN_EN;

