------------------------------------------------------------------------------
--  This file is a part of the GRLIB VHDL IP LIBRARY
--  Copyright (C) 2015, Cobham Gaisler AB - all rights reserved.
--
-- ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN 
-- ACCORDANCE WITH THE GAISLER LICENSE AGREEMENT AND MUST BE APPROVED 
-- IN ADVANCE IN WRITING. 
-----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.all;

entity grlfpw_0_unisim is
port(
  rst :  in std_logic;
  clk :  in std_logic;
  holdn :  in std_logic;
  cpi_flush :  in std_logic;
  cpi_exack :  in std_logic;
  cpi_a_rs1 : in std_logic_vector(4 downto 0);
  cpi_d_pc : in std_logic_vector(31 downto 0);
  cpi_d_inst : in std_logic_vector(31 downto 0);
  cpi_d_cnt : in std_logic_vector(1 downto 0);
  cpi_d_trap :  in std_logic;
  cpi_d_annul :  in std_logic;
  cpi_d_pv :  in std_logic;
  cpi_a_pc : in std_logic_vector(31 downto 0);
  cpi_a_inst : in std_logic_vector(31 downto 0);
  cpi_a_cnt : in std_logic_vector(1 downto 0);
  cpi_a_trap :  in std_logic;
  cpi_a_annul :  in std_logic;
  cpi_a_pv :  in std_logic;
  cpi_e_pc : in std_logic_vector(31 downto 0);
  cpi_e_inst : in std_logic_vector(31 downto 0);
  cpi_e_cnt : in std_logic_vector(1 downto 0);
  cpi_e_trap :  in std_logic;
  cpi_e_annul :  in std_logic;
  cpi_e_pv :  in std_logic;
  cpi_m_pc : in std_logic_vector(31 downto 0);
  cpi_m_inst : in std_logic_vector(31 downto 0);
  cpi_m_cnt : in std_logic_vector(1 downto 0);
  cpi_m_trap :  in std_logic;
  cpi_m_annul :  in std_logic;
  cpi_m_pv :  in std_logic;
  cpi_x_pc : in std_logic_vector(31 downto 0);
  cpi_x_inst : in std_logic_vector(31 downto 0);
  cpi_x_cnt : in std_logic_vector(1 downto 0);
  cpi_x_trap :  in std_logic;
  cpi_x_annul :  in std_logic;
  cpi_x_pv :  in std_logic;
  cpi_lddata : in std_logic_vector(31 downto 0);
  cpi_dbg_enable :  in std_logic;
  cpi_dbg_write :  in std_logic;
  cpi_dbg_fsr :  in std_logic;
  cpi_dbg_addr : in std_logic_vector(4 downto 0);
  cpi_dbg_data : in std_logic_vector(31 downto 0);
  cpo_data : out std_logic_vector(31 downto 0);
  cpo_exc :  out std_logic;
  cpo_cc : out std_logic_vector(1 downto 0);
  cpo_ccv :  out std_logic;
  cpo_ldlock :  out std_logic;
  cpo_holdn :  out std_logic;
  cpo_dbg_data : out std_logic_vector(31 downto 0);
  rfi1_rd1addr : out std_logic_vector(3 downto 0);
  rfi1_rd2addr : out std_logic_vector(3 downto 0);
  rfi1_wraddr : out std_logic_vector(3 downto 0);
  rfi1_wrdata : out std_logic_vector(31 downto 0);
  rfi1_ren1 :  out std_logic;
  rfi1_ren2 :  out std_logic;
  rfi1_wren :  out std_logic;
  rfi2_rd1addr : out std_logic_vector(3 downto 0);
  rfi2_rd2addr : out std_logic_vector(3 downto 0);
  rfi2_wraddr : out std_logic_vector(3 downto 0);
  rfi2_wrdata : out std_logic_vector(31 downto 0);
  rfi2_ren1 :  out std_logic;
  rfi2_ren2 :  out std_logic;
  rfi2_wren :  out std_logic;
  rfo1_data1 : in std_logic_vector(31 downto 0);
  rfo1_data2 : in std_logic_vector(31 downto 0);
  rfo2_data1 : in std_logic_vector(31 downto 0);
  rfo2_data2 : in std_logic_vector(31 downto 0));
end grlfpw_0_unisim;

architecture beh of grlfpw_0_unisim is
  signal \GRLFPC20.R.FSR.RD\ : std_logic_vector(1 downto 0);
  signal \GRLFPC20.FPO.EXC\ : std_logic_vector(3 downto 1);
  signal \GRLFPC20.R.STATE\ : std_logic_vector(1 downto 0);
  signal \GRLFPC20.R.I.INST\ : std_logic_vector(31 downto 0);
  signal \GRLFPC20.R.FSR.TEM\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.R.I.EXC\ : std_logic_vector(5 downto 0);
  signal \GRLFPC20.R.FSR.AEXC\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.R.A.RS1\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.R.A.RS2\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.R.I.PC\ : std_logic_vector(31 downto 2);
  signal \GRLFPC20.R.FSR.CEXC\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.R.FSR.FTT\ : std_logic_vector(2 downto 0);
  signal \GRLFPC20.R.I.CC\ : std_logic_vector(1 downto 0);
  signal \GRLFPC20.R.I.RES\ : std_logic_vector(63 downto 0);
  signal \GRLFPC20.COMB.V.I.RES_1\ : std_logic_vector(63 downto 29);
  signal \GRLFPC20.COMB.V.FSR.FTT_1\ : std_logic_vector(2 downto 0);
  signal \GRLFPC20.R.A.RF1REN\ : std_logic_vector(2 downto 1);
  signal \GRLFPC20.R.A.RF2REN\ : std_logic_vector(2 downto 1);
  signal \GRLFPC20.COMB.V.FSR.FCC_1\ : std_logic_vector(1 downto 0);
  signal \GRLFPC20.COMB.V.FSR.AEXC_1\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.COMB.V.FSR.CEXC_1\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.COMB.V.FSR.TEM_1\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.COMB.V.E.STDATA_1\ : std_logic_vector(31 downto 0);
  signal \GRLFPC20.COMB.RS1_1\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\ : std_logic_vector(16 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_25\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_DIVMULTV\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\ : std_logic_vector(85 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\ : std_logic_vector(377 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.MIXOIN\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\ : std_logic_vector(57 downto 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\ : std_logic_vector(113 downto 58);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\ : std_logic_vector(53 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN17_XZXBUS\ : std_logic_vector(1 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\ : std_logic_vector(11 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14\ : std_logic_vector(77 to 77);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_18\ : std_logic_vector(74 to 74);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_21\ : std_logic_vector(40 to 40);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_49\ : std_logic_vector(258 to 258);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_10\ : std_logic_vector(10 to 10);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\ : std_logic_vector(375 downto 58);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_13\ : std_logic_vector(3 to 3);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_14\ : std_logic_vector(4 to 4);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\ : std_logic_vector(9 downto 7);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1\ : std_logic_vector(7 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_61\ : std_logic_vector(52 to 52);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.SI_118\ : std_logic_vector(51 to 51);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\ : std_logic_vector(57 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\ : std_logic_vector(62 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRLOI\ : std_logic_vector(34 downto 29);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\ : std_logic_vector(57 downto 2);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\ : std_logic_vector(57 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN8_TEMP\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\ : std_logic_vector(57 downto 2);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\ : std_logic_vector(9 downto 4);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\ : std_logic_vector(18 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_DATA_TMP\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.COMB.V.STATE_1\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.COMB.V.FSR.RD_1\ : std_logic_vector(1 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_50\ : std_logic_vector(316 to 316);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\ : std_logic_vector(54 downto 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\ : std_logic_vector(55 downto 10);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\ : std_logic_vector(54 downto 3);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\ : std_logic_vector(1 to 1);
  signal \GRLFPC20.COMB.WRDATA_4\ : std_logic_vector(62 downto 0);
  signal \GRLFPC20.FPI.OP2\ : std_logic_vector(62 downto 32);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\ : std_logic_vector(57 downto 33);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\ : std_logic_vector(83 downto 61);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\ : std_logic_vector(53 downto 51);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\ : std_logic_vector(57 downto 19);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_114\ : std_logic_vector(56 to 56);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M12\ : std_logic_vector(2 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M13\ : std_logic_vector(2 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M8\ : std_logic_vector(2 downto 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2\ : std_logic_vector(3 to 3);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14_2\ : std_logic_vector(77 to 77);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_11\ : std_logic_vector(7 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_10\ : std_logic_vector(7 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\ : std_logic_vector(7 downto 3);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SALSBS_2\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\ : std_logic_vector(8 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\ : std_logic_vector(2 to 2);
  signal \GRLFPC20.FPI.OP1\ : std_logic_vector(62 downto 32);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SALSBS_1\ : std_logic_vector(1 to 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_9\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_19\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\ : std_logic_vector(67 to 67);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\ : std_logic_vector(57 downto 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS_2\ : std_logic_vector(1 to 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\ : std_logic_vector(3 to 3);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_WQSTSETS\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\ : std_logic_vector(56 downto 33);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.U_RDN_1\ : std_logic_vector(1 to 1);
  signal \GRLFPC20.COMB.V.STATE_9\ : std_logic_vector(1 downto 0);
  signal \GRLFPC20.COMB.V.A.RF2REN_1\ : std_logic_vector(2 downto 1);
  signal \GRLFPC20.COMB.V.A.RF1REN_1\ : std_logic_vector(1 to 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SBLSBS_2\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.R.I.EXC_M\ : std_logic_vector(2 to 2);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_2\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_S0\ : std_logic_vector(3 to 3);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_T_3\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_14\ : std_logic_vector(172 downto 141);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41\ : std_logic_vector(254 downto 253);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.LIB\ : std_logic_vector(1 to 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.RESULT\ : std_logic_vector(2 to 2);
  signal \GRLFPC20.COMB.V.FSR.FCC_1_M0\ : std_logic_vector(1 downto 0);
  signal \GRLFPC20.COMB.V.FSR.AEXC_1_M0\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.FPO.EXP\ : std_logic_vector(10 downto 0);
  signal \GRLFPC20.FPO.FRAC\ : std_logic_vector(54 downto 3);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.SI_64\ : std_logic_vector(49 to 49);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.SI_6\ : std_logic_vector(51 to 51);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.SI_63\ : std_logic_vector(50 to 50);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.SI_120\ : std_logic_vector(49 to 49);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_5\ : std_logic_vector(52 to 52);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.SI_119\ : std_logic_vector(50 to 50);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.SI_79\ : std_logic_vector(34 to 34);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.SI_21\ : std_logic_vector(36 to 36);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.SI_78\ : std_logic_vector(35 to 35);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.SI_134\ : std_logic_vector(35 to 35);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.SI_19\ : std_logic_vector(38 to 38);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.SI_133\ : std_logic_vector(36 to 36);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.SI_18\ : std_logic_vector(39 to 39);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.SI_74\ : std_logic_vector(39 to 39);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.SI_16\ : std_logic_vector(41 to 41);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.SI_130\ : std_logic_vector(39 to 39);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.SI_15\ : std_logic_vector(42 to 42);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.SI_72\ : std_logic_vector(41 to 41);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.SI_14\ : std_logic_vector(43 to 43);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.SI_71\ : std_logic_vector(42 to 42);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.SI_70\ : std_logic_vector(43 to 43);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.SI_127\ : std_logic_vector(42 to 42);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.SI_12\ : std_logic_vector(45 to 45);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.SI_126\ : std_logic_vector(43 to 43);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.SI_11\ : std_logic_vector(46 to 46);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.SI_68\ : std_logic_vector(45 to 45);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.SI_125\ : std_logic_vector(44 to 44);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.SI_10\ : std_logic_vector(47 to 47);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.SI_124\ : std_logic_vector(45 to 45);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.SI_9\ : std_logic_vector(48 to 48);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.SI_8\ : std_logic_vector(49 to 49);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.SI_65\ : std_logic_vector(48 to 48);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.SI_37\ : std_logic_vector(20 to 20);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.SI_36\ : std_logic_vector(21 to 21);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.SI_93\ : std_logic_vector(20 to 20);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.SI_149\ : std_logic_vector(20 to 20);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.SI_34\ : std_logic_vector(23 to 23);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.SI_33\ : std_logic_vector(24 to 24);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.SI_32\ : std_logic_vector(25 to 25);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.SI_30\ : std_logic_vector(27 to 27);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.SI_87\ : std_logic_vector(26 to 26);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.SI_29\ : std_logic_vector(28 to 28);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.SI_28\ : std_logic_vector(29 to 29);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.SI_85\ : std_logic_vector(28 to 28);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.SI_84\ : std_logic_vector(29 to 29);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.SI_26\ : std_logic_vector(31 to 31);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.SI_140\ : std_logic_vector(29 to 29);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.SI_25\ : std_logic_vector(32 to 32);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.SI_139\ : std_logic_vector(30 to 30);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.SI_24\ : std_logic_vector(33 to 33);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.SI_23\ : std_logic_vector(34 to 34);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.SI_80\ : std_logic_vector(33 to 33);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.SI_103\ : std_logic_vector(10 to 10);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.SI_160\ : std_logic_vector(9 to 9);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.SI_45\ : std_logic_vector(12 to 12);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.SI_44\ : std_logic_vector(13 to 13);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.SI_101\ : std_logic_vector(12 to 12);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.SI_43\ : std_logic_vector(14 to 14);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.SI_100\ : std_logic_vector(13 to 13);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.SI_41\ : std_logic_vector(16 to 16);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.SI_98\ : std_logic_vector(15 to 15);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.SI_155\ : std_logic_vector(14 to 14);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.SI_40\ : std_logic_vector(17 to 17);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.SI_97\ : std_logic_vector(16 to 16);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.SI_154\ : std_logic_vector(15 to 15);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.SI_39\ : std_logic_vector(18 to 18);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.SI_38\ : std_logic_vector(19 to 19);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.SI_95\ : std_logic_vector(18 to 18);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.SI_152\ : std_logic_vector(17 to 17);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.SI_167\ : std_logic_vector(2 to 2);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.SI_51\ : std_logic_vector(6 to 6);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.SI_108\ : std_logic_vector(5 to 5);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.SI_165\ : std_logic_vector(4 to 4);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.SI_50\ : std_logic_vector(7 to 7);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.SI_106\ : std_logic_vector(7 to 7);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.SI_163\ : std_logic_vector(6 to 6);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.SI_48\ : std_logic_vector(9 to 9);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.SI_105\ : std_logic_vector(8 to 8);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.SI_47\ : std_logic_vector(10 to 10);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SBLSBS_1\ : std_logic_vector(1 to 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.SI_56\ : std_logic_vector(1 to 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_113\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SCLSBS_1\ : std_logic_vector(1 to 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.SI_55\ : std_logic_vector(2 to 2);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.SI_112\ : std_logic_vector(1 to 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.SI_54\ : std_logic_vector(3 to 3);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\ : std_logic_vector(12 downto 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_I\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9\ : std_logic_vector(58 downto 27);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3\ : std_logic_vector(55 downto 6);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_16_TZ\ : std_logic_vector(54 to 54);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_21_0_1_TZ\ : std_logic_vector(40 to 40);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_13\ : std_logic_vector(11 to 11);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\ : std_logic_vector(62 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_7_TZ\ : std_logic_vector(56 to 56);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_16_0\ : std_logic_vector(52 to 52);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_15_1\ : std_logic_vector(36 to 36);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_17_0\ : std_logic_vector(11 to 11);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_7_1\ : std_logic_vector(25 to 25);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_5_0\ : std_logic_vector(48 to 48);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_23_0\ : std_logic_vector(47 to 47);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_8_0\ : std_logic_vector(54 to 54);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A26_22_0\ : std_logic_vector(60 to 60);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_10_1\ : std_logic_vector(61 to 61);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_0\ : std_logic_vector(15 downto 11);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_9_0\ : std_logic_vector(47 to 47);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_1_0\ : std_logic_vector(36 to 36);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_2_0\ : std_logic_vector(5 to 5);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A12_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0_0_A2_0\ : std_logic_vector(0 to 0);
  signal CPI_D_INST_I : std_logic_vector(6 to 6);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_I\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_25_I\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\ : std_logic_vector(69 downto 42);
  signal \GRLFPC20.COMB.V.STATE_1_IV_I\ : std_logic_vector(1 to 1);
  signal \GRLFPC20.RS1_1_0_0\ : std_logic_vector(4 downto 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1_0\ : std_logic_vector(5 downto 4);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1_2\ : std_logic_vector(6 to 6);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1_3\ : std_logic_vector(6 to 6);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A22_2_0\ : std_logic_vector(53 to 53);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_7_0\ : std_logic_vector(4 to 4);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_22_0\ : std_logic_vector(54 to 54);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A24_0\ : std_logic_vector(59 to 59);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A22_16_0\ : std_logic_vector(53 to 53);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A30_14_0\ : std_logic_vector(58 to 58);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_20_0\ : std_logic_vector(57 to 57);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_6_1\ : std_logic_vector(25 to 25);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_7_0\ : std_logic_vector(48 to 48);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A30_10_1\ : std_logic_vector(58 to 58);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_3_1\ : std_logic_vector(32 to 32);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A24_7_0\ : std_logic_vector(59 to 59);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_11_0\ : std_logic_vector(19 to 19);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A26_3_1\ : std_logic_vector(60 to 60);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_I_A2_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_I_A2_1\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_I_A2_2\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_I_A2_3\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_I_A2_4\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A24_10_1\ : std_logic_vector(59 to 59);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_9_1\ : std_logic_vector(57 to 57);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A24_19_1\ : std_logic_vector(59 to 59);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A30_23_0\ : std_logic_vector(58 to 58);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_0\ : std_logic_vector(4 to 4);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A30_4_0\ : std_logic_vector(58 to 58);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A30_4_1\ : std_logic_vector(58 to 58);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_6_0\ : std_logic_vector(57 to 57);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_1_1\ : std_logic_vector(36 downto 7);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_0_0\ : std_logic_vector(25 to 25);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_9_0\ : std_logic_vector(55 to 55);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A12_0_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_9_0\ : std_logic_vector(25 to 25);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_2_0\ : std_logic_vector(52 to 52);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_6_0\ : std_logic_vector(52 to 52);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_8_1\ : std_logic_vector(13 to 13);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_8_1\ : std_logic_vector(19 to 19);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_3_2\ : std_logic_vector(19 to 19);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_9_1\ : std_logic_vector(52 to 52);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_1_1\ : std_logic_vector(32 to 32);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_6_1\ : std_logic_vector(32 to 32);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_7_0\ : std_logic_vector(52 to 52);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.EXTEND.TEMP_0\ : std_logic_vector(1 to 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A8_5_2\ : std_logic_vector(62 to 62);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_11_0\ : std_logic_vector(52 to 52);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_2_A2_0_A2_0\ : std_logic_vector(51 to 51);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A22_11_0\ : std_logic_vector(53 to 53);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_0_0\ : std_logic_vector(6 to 6);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_6_0\ : std_logic_vector(47 to 47);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_0_A2_0_A2_0\ : std_logic_vector(51 to 51);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0\ : std_logic_vector(50 downto 14);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1\ : std_logic_vector(50 downto 5);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\ : std_logic_vector(62 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\ : std_logic_vector(61 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2\ : std_logic_vector(61 downto 3);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_0\ : std_logic_vector(61 downto 24);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5\ : std_logic_vector(61 downto 13);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_1\ : std_logic_vector(18 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0\ : std_logic_vector(59 downto 18);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\ : std_logic_vector(59 downto 6);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_O2_0\ : std_logic_vector(24 to 24);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_1\ : std_logic_vector(49 downto 5);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0_0\ : std_logic_vector(35 to 35);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15_0_0\ : std_logic_vector(16 to 16);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15_1\ : std_logic_vector(16 to 16);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_1\ : std_logic_vector(36 downto 6);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0\ : std_logic_vector(59 downto 6);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0\ : std_logic_vector(59 downto 6);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8\ : std_logic_vector(58 downto 19);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_0\ : std_logic_vector(54 downto 6);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_0\ : std_logic_vector(59 downto 27);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7\ : std_logic_vector(59 downto 6);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4\ : std_logic_vector(59 downto 6);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_1\ : std_logic_vector(58 downto 13);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2\ : std_logic_vector(50 downto 4);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_0\ : std_logic_vector(51 downto 4);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_0\ : std_logic_vector(51 downto 4);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_0\ : std_logic_vector(51 downto 4);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_3\ : std_logic_vector(4 to 4);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3\ : std_logic_vector(50 downto 5);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_4\ : std_logic_vector(5 to 5);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_1\ : std_logic_vector(58 downto 6);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_1\ : std_logic_vector(57 downto 19);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_1\ : std_logic_vector(59 to 59);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_0\ : std_logic_vector(60 downto 11);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_4\ : std_logic_vector(60 downto 47);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_5\ : std_logic_vector(60 downto 47);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_7\ : std_logic_vector(60 downto 11);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_0_0\ : std_logic_vector(47 to 47);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_1_0\ : std_logic_vector(60 downto 47);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2_0\ : std_logic_vector(60 downto 47);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_3_0\ : std_logic_vector(47 downto 11);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_4_0\ : std_logic_vector(56 downto 11);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_5_0\ : std_logic_vector(47 downto 11);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_6_0\ : std_logic_vector(56 downto 47);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_6_1\ : std_logic_vector(47 to 47);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2_1\ : std_logic_vector(60 downto 11);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2\ : std_logic_vector(56 downto 11);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_3\ : std_logic_vector(60 downto 11);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_6\ : std_logic_vector(56 downto 11);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_7_0\ : std_logic_vector(56 downto 11);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_1_1\ : std_logic_vector(11 to 11);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_1\ : std_logic_vector(57 to 57);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_11\ : std_logic_vector(57 downto 52);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_13\ : std_logic_vector(57 to 57);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_0\ : std_logic_vector(31 to 31);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_2\ : std_logic_vector(31 to 31);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_5\ : std_logic_vector(31 to 31);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_0_0\ : std_logic_vector(31 to 31);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_1_0\ : std_logic_vector(31 to 31);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_2_0\ : std_logic_vector(31 to 31);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_3_0\ : std_logic_vector(31 to 31);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_4_1\ : std_logic_vector(31 to 31);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_5_1\ : std_logic_vector(31 to 31);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_6_0\ : std_logic_vector(31 to 31);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_6_1\ : std_logic_vector(31 to 31);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_7_0\ : std_logic_vector(31 to 31);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_0_1\ : std_logic_vector(31 to 31);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7_0\ : std_logic_vector(33 downto 19);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7_1\ : std_logic_vector(58 downto 52);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8_2\ : std_logic_vector(58 to 58);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8_0\ : std_logic_vector(54 to 54);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8_1\ : std_logic_vector(54 to 54);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9_0\ : std_logic_vector(54 to 54);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_12\ : std_logic_vector(54 to 54);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_0_1\ : std_logic_vector(60 to 60);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_5_1\ : std_logic_vector(60 to 60);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_6_2\ : std_logic_vector(60 to 60);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2_2\ : std_logic_vector(60 to 60);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_1\ : std_logic_vector(49 to 49);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_2\ : std_logic_vector(49 to 49);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_2\ : std_logic_vector(49 to 49);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_1\ : std_logic_vector(56 to 56);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_8\ : std_logic_vector(56 to 56);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_4_1\ : std_logic_vector(51 to 51);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_5_0\ : std_logic_vector(51 to 51);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_5_1\ : std_logic_vector(51 to 51);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_1\ : std_logic_vector(51 to 51);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0_0_O2_0\ : std_logic_vector(2 to 2);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0_0_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.COMB.V.FSR.CEXC_1_IV_1\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.COMB.V.FSR.CEXC_1_IV_0\ : std_logic_vector(2 to 2);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8_1\ : std_logic_vector(57 to 57);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8_0_0\ : std_logic_vector(57 to 57);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8_1_1\ : std_logic_vector(57 to 57);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_1_1\ : std_logic_vector(28 downto 20);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.RESULT_IV_0\ : std_logic_vector(1 to 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_26_A0_1\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_1\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_28_0\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.R.X.RDD_TMP_D_ARRAY_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.R.X.SEQERR_TMP_D_ARRAY_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\ : std_logic_vector(30 downto 8);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_FAST\ : std_logic_vector(19 downto 8);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_REP1\ : std_logic_vector(17 downto 16);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_REP2\ : std_logic_vector(17 downto 16);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST\ : std_logic_vector(376 downto 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_FAST\ : std_logic_vector(374 to 374);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_FAST\ : std_logic_vector(17 downto 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_DIVMULTV_FAST\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_REP1\ : std_logic_vector(9 downto 3);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_FAST\ : std_logic_vector(10 to 10);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\ : std_logic_vector(236 downto 232);
  signal \GRLFPC20.COMB.V.A.RF1REN_1_0\ : std_logic_vector(2 to 2);
  signal \GRLFPC20.COMB.RS1_1_0_0\ : std_logic_vector(4 downto 1);
  signal \GRLFPC20.COMB.RS2_1_0\ : std_logic_vector(4 downto 1);
  signal \GRLFPC20.COMB.RS2_1DUP\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_2_0_E\ : std_logic_vector(65 to 65);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_E_0_E\ : std_logic_vector(69 to 69);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_5_0_E\ : std_logic_vector(1 to 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_4_0_E\ : std_logic_vector(2 to 2);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_6_0_E\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14_0_E\ : std_logic_vector(77 to 77);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_16_0_E\ : std_logic_vector(6 to 6);
  signal \GRLFPC20.COMB.V.STATE_9_I\ : std_logic_vector(0 to 0);
  signal CPO_EXC_1 : std_logic ;
  signal NN_1 : std_logic ;
  signal CPO_CC_3 : std_logic ;
  signal NN_2 : std_logic ;
  signal NN_3 : std_logic ;
  signal \GRLFPC20.FPI.START\ : std_logic ;
  signal \GRLFPC20.R.I.EXEC\ : std_logic ;
  signal \GRLFPC20.R.MK.BUSY\ : std_logic ;
  signal \GRLFPC20.R.X.LD\ : std_logic ;
  signal \GRLFPC20.R.X.AFSR\ : std_logic ;
  signal \GRLFPC20.R.X.SEQERR\ : std_logic ;
  signal \GRLFPC20.R.X.FPOP\ : std_logic ;
  signal \GRLFPC20.R.A.RS1D\ : std_logic ;
  signal \GRLFPC20.R.A.RS2D\ : std_logic ;
  signal \GRLFPC20.R.A.AFQ\ : std_logic ;
  signal \GRLFPC20.R.MK.RST\ : std_logic ;
  signal \GRLFPC20.R.MK.RST2\ : std_logic ;
  signal \GRLFPC20.R.MK.HOLDN1\ : std_logic ;
  signal \GRLFPC20.R.E.FPOP\ : std_logic ;
  signal \GRLFPC20.R.M.FPOP\ : std_logic ;
  signal \GRLFPC20.R.A.ST\ : std_logic ;
  signal \GRLFPC20.R.A.AFSR\ : std_logic ;
  signal \GRLFPC20.R.MK.HOLDN2\ : std_logic ;
  signal \GRLFPC20.R.I.V\ : std_logic ;
  signal \GRLFPC20.R.M.LD\ : std_logic ;
  signal \GRLFPC20.R.E.LD\ : std_logic ;
  signal \GRLFPC20.R.A.LD\ : std_logic ;
  signal \GRLFPC20.R.A.FPOP\ : std_logic ;
  signal \GRLFPC20.R.MK.LDOP\ : std_logic ;
  signal \GRLFPC20.COMB.V.X.AFQ_1\ : std_logic ;
  signal \GRLFPC20.R.M.AFQ\ : std_logic ;
  signal \GRLFPC20.COMB.V.X.AFSR_1\ : std_logic ;
  signal \GRLFPC20.R.M.AFSR\ : std_logic ;
  signal \GRLFPC20.COMB.V.X.FPOP_1\ : std_logic ;
  signal \GRLFPC20.COMB.V.X.LD_1\ : std_logic ;
  signal \GRLFPC20.COMB.V.M.AFQ_1\ : std_logic ;
  signal \GRLFPC20.R.E.AFQ\ : std_logic ;
  signal \GRLFPC20.COMB.V.M.AFSR_1\ : std_logic ;
  signal \GRLFPC20.R.E.AFSR\ : std_logic ;
  signal \GRLFPC20.COMB.V.M.FPOP_1\ : std_logic ;
  signal \GRLFPC20.COMB.V.M.LD_1\ : std_logic ;
  signal \GRLFPC20.COMB.V.E.AFQ_1\ : std_logic ;
  signal \GRLFPC20.COMB.V.E.AFSR_1\ : std_logic ;
  signal \GRLFPC20.N_2931_1\ : std_logic ;
  signal \GRLFPC20.COMB.V.E.LD_1\ : std_logic ;
  signal \GRLFPC20.R.X.AFQ\ : std_logic ;
  signal \GRLFPC20.R.A.MOV\ : std_logic ;
  signal \GRLFPC20.R.I.RDD\ : std_logic ;
  signal \GRLFPC20.R.X.RDD\ : std_logic ;
  signal \GRLFPC20.R.MK.BUSY2\ : std_logic ;
  signal \GRLFPC20.R.FSR.NONSTD\ : std_logic ;
  signal \GRLFPC20.COMB.V.MK.BUSY2_2\ : std_logic ;
  signal \GRLFPC20.COMB.V.MK.RST_1\ : std_logic ;
  signal \GRLFPC20.COMB.V.MK.BUSY_2\ : std_logic ;
  signal \GRLFPC20.V.I.V_3_SQMUXA\ : std_logic ;
  signal \GRLFPC20.N_1858\ : std_logic ;
  signal \GRLFPC20.N_2102\ : std_logic ;
  signal \GRLFPC20.N_1338\ : std_logic ;
  signal \GRLFPC20.COMB.V.FSR.AEXC_1_SN.N_7_MUX\ : std_logic ;
  signal \GRLFPC20.COMB.V.FSR.NONSTD_1\ : std_logic ;
  signal \GRLFPC20.N_1704\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN3_NOTRESETORUNIMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9252\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9260\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_11\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_18\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_25\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_32\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_39\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_53\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_60\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_67\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_81\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_88\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_95\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_102\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_109\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_116\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_123\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_130\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_N_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_N_11\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_N_18\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_N_25\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12030\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12045\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN2_NOTDECODEDUNIMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_453\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_457\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_499\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_513\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_515\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_519\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_521\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_523\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_537\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_541\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_544\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_548\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_550\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_552\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_554\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_559\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_753\ : std_logic ;
  signal \GRLFPC20.COMB.RS2D_1\ : std_logic ;
  signal \GRLFPC20.COMB.RS1D_1\ : std_logic ;
  signal \GRLFPC20.COMB.V.A.AFQ_1\ : std_logic ;
  signal \GRLFPC20.COMB.V.A.SEQERR_1\ : std_logic ;
  signal \GRLFPC20.COMB.V.A.AFSR_1\ : std_logic ;
  signal \GRLFPC20.COMB.V.A.ST_1\ : std_logic ;
  signal \GRLFPC20.N_1312\ : std_logic ;
  signal \GRLFPC20.COMB.V.A.LD_1\ : std_logic ;
  signal \GRLFPC20.COMB.RDD_1\ : std_logic ;
  signal \GRLFPC20.N_865\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9144\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9084\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_4_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\ : std_logic ;
  signal \GRLFPC20.FPI.LDOP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8654\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7944\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7936\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7884\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7708\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_187\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9154\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9094\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8646\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8641\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8636\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7931\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7926\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7876\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7700\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7871\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7695\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7866\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7690\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8223\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_601\ : std_logic ;
  signal \GRLFPC20.WRADDR_0_SQMUXA\ : std_logic ;
  signal \GRLFPC20.N_1562\ : std_logic ;
  signal \GRLFPC20.COMB.RDD_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SS0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10948_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_143\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9670_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_125\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10824_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2454_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_369\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_222\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9700_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10895\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10661\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9861_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_304\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1661\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1971\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1562\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2701\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2669\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2630\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2605\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9389_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9666_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9666_1_I_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9461_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_717\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9738_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_783\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1019_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9790_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_406\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9863_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10224\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9394_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_715\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9850_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9667_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10207_I_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_795\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10211\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9549_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_746\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_831\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10025_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_749\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_909\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9577\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2601\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1335\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_777\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2590\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1192\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1232\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2721\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1272\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_157_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1344\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_742\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_921\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2337\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_291_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9176\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9067\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9127\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9116\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_4_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8364\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7977\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8687\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8366\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8358\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7741\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8362\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9249\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12250\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9316\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9330_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9324_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9296_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9326\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9858_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9320_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9975_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_747_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9323\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9321_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9604_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9671_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9652_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9797_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_52\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10734\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9314\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9492_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9338\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9338_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_990_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_59\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9973_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9328\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9972_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1230\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_720\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9657_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_328\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12132\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9558_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9318\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9993\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9610_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9390_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10531\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9969_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_261\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10869\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9968_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_782\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1776\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1169\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_722\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_SM12\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_SS0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8535\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8533\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_584\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8532\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12036\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8551\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8550\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8549\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8548\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8546\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8545\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_93\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1323\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1137\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12041\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12032\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8547\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8534\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_SS9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12249\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2505_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2150\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2800\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_776\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2635\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2583\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_775\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9561\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9600_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9551_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1725\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2448\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_11378\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2724\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2584\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2591\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_766\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2230\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2156\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2151\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1654\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10088\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2831\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_134_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_234\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2606\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9506_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2594\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_202\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9925_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9655_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9404_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_759\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1650\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1336\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2602\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1234\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_741\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2608\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1170\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_789\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1133\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1025\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2206\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1592\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_982\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_989\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_966\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9785_1_I_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1132_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12131\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2600\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1229\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_995_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2730\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10146\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9503_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10157\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10158\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10157_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10456\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2400\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.OPREXCSHFT.UN3_OPREXC\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2216\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1536_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2255\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1653\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_534\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2233\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_765\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_135\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2758\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2140\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2762\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9663\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_85\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2166\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1283\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9453_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1282\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2764\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2403\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1039\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1149\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_906\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10410\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_732\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_751_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1331\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9508_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_0_SN_N_7_MUX\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_0_SN_N_6_MUX\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1710\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1648\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2445\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2229_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1711\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2159\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2447\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2475\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10654\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9605_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8114\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2842\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2774\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_907\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10626_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10892\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10929\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10917\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10927_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10926\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10640\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10925\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.MIFROMINST\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.TEMP_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_981\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_979\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_978\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_965\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_289\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1333\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CONDMUXMULXFF.UN5_NOTSQRTLFTCC\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7498_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO0_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9169\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9139\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9109\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9079\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_812_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_811_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO1_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN18_GEN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN12_GEN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN10_NOTPROP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.NOTPROP_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.NOTPROP_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN1_NOTPROP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.STKGEN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN16_NOTPROP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN22_NOTPROP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN20_STKOUT\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.STKGEN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9969_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10164\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10884\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10882\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10767_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10888_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9994_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9555_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9505_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9665_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10893\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10891\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10891_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10891_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_76\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10693_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10163\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10167\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7596\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8109\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN1_S_14\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.ENTRYPOINT\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2695\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9563_1\ : std_logic ;
  signal \GRLFPC20.N_878\ : std_logic ;
  signal \GRLFPC20.COMB.FPDECODE.RS1D5\ : std_logic ;
  signal \GRLFPC20.N_940\ : std_logic ;
  signal \GRLFPC20.N_3128\ : std_logic ;
  signal \GRLFPC20.N_3129\ : std_logic ;
  signal \GRLFPC20.N_3127\ : std_logic ;
  signal \GRLFPC20.N_3123\ : std_logic ;
  signal \GRLFPC20.COMB.RDD_1.I9_MUX\ : std_logic ;
  signal \GRLFPC20.RS1D_CNST.N_7\ : std_logic ;
  signal \GRLFPC20.COMB.LOCKGEN.LOCKI\ : std_logic ;
  signal \GRLFPC20.COMB.RS1V_1\ : std_logic ;
  signal \GRLFPC20.RS1D_CNST\ : std_logic ;
  signal \GRLFPC20.N_3074\ : std_logic ;
  signal \GRLFPC20.N_3116\ : std_logic ;
  signal \GRLFPC20.N_3117\ : std_logic ;
  signal \GRLFPC20.N_3084\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN10_S_MOV\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9913_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2517_2\ : std_logic ;
  signal \GRLFPC20.N_3106\ : std_logic ;
  signal \GRLFPC20.N_3079\ : std_logic ;
  signal \GRLFPC20.N_3120\ : std_logic ;
  signal \GRLFPC20.N_3083_1\ : std_logic ;
  signal \GRLFPC20.N_925\ : std_logic ;
  signal \GRLFPC20.N_3081\ : std_logic ;
  signal \GRLFPC20.N_2962\ : std_logic ;
  signal \GRLFPC20.RS1V_0_SQMUXA_1\ : std_logic ;
  signal \GRLFPC20.N_1583\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN3_NOTAZERODENORM\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8581\ : std_logic ;
  signal \GRLFPC20.V.I.EXEC_0_SQMUXA\ : std_logic ;
  signal \GRLFPC20.N_1528\ : std_logic ;
  signal \GRLFPC20.R.X.SEQERR_M\ : std_logic ;
  signal \GRLFPC20.N_1494\ : std_logic ;
  signal \GRLFPC20.WREN1_1_SQMUXA\ : std_logic ;
  signal \GRLFPC20.COMB.WREN1_2_M\ : std_logic ;
  signal \GRLFPC20.N_1475\ : std_logic ;
  signal \GRLFPC20.N_2015\ : std_logic ;
  signal \GRLFPC20.N_1295\ : std_logic ;
  signal \GRLFPC20.COMB.UN1_ANNULFPU\ : std_logic ;
  signal \GRLFPC20.N_2395\ : std_logic ;
  signal \GRLFPC20.COMB.V.E.STDATA2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\ : std_logic ;
  signal \GRLFPC20.N_2112\ : std_logic ;
  signal \GRLFPC20.N_2045\ : std_logic ;
  signal \GRLFPC20.N_1317\ : std_logic ;
  signal \GRLFPC20.COMB.FPDECODE.ST\ : std_logic ;
  signal \GRLFPC20.RS1V_0_SQMUXA\ : std_logic ;
  signal \GRLFPC20.COMB.UN1_FPCI_4\ : std_logic ;
  signal \GRLFPC20.COMB.UN1_R.A.RS1_1\ : std_logic ;
  signal \GRLFPC20.N_3109\ : std_logic ;
  signal \GRLFPC20.N_2512\ : std_logic ;
  signal \GRLFPC20.COMB.V.A.AFQ_1_1\ : std_logic ;
  signal \GRLFPC20.N_1138\ : std_logic ;
  signal \GRLFPC20.N_1142\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.NOTABORTWB\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8306\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8212\ : std_logic ;
  signal \GRLFPC20.N_3050\ : std_logic ;
  signal \GRLFPC20.N_2000\ : std_logic ;
  signal \GRLFPC20.N_2397\ : std_logic ;
  signal \GRLFPC20.N_2388\ : std_logic ;
  signal \GRLFPC20.V.STATE_2_SQMUXA\ : std_logic ;
  signal \GRLFPC20.N_1421\ : std_logic ;
  signal \GRLFPC20.N_2385\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8284\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9099\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9159\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9163\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9103\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8580\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.UN84_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8539\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8658\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7948\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7888\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7712\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9167\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9165\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9107\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9105\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7894\ : std_logic ;
  signal \GRLFPC20.N_2103\ : std_logic ;
  signal \GRLFPC20.COMB.ANNULRES_1\ : std_logic ;
  signal \GRLFPC20.COMB.V.I.EXEC_5\ : std_logic ;
  signal \GRLFPC20.N_1597\ : std_logic ;
  signal \GRLFPC20.COMB.UN15_HOLDN\ : std_logic ;
  signal \GRLFPC20.FPO.SIGN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9257\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SFTLFT.AREGXORBREG\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8230\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8218\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8235\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8233\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8231\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8232\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8228\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8244\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8243\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8241\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8237\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8215\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8211\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8246\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8238\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8236\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8227\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8219\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8213\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8214\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8209\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8210\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8208\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8207\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8205\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8201\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8199\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8200\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8198\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1086\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8245\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8234\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8202\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8203\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8204\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8206\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8690\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7979\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12044\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7512\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO0_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO2_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO0_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO0_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8686\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8685\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7976\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7740\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_58_2.CO1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.UN348_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7975\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7739\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_2.CO3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_2.CO2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.UN3_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8815\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8830\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8822\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8825\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8821\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8814\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8807\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8810\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9922_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12195\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_409\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1553_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10016\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10035\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10006\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10030_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_768_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10024\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10023\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10022\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9971\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9161\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9101\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9158\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9098\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8292\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8321\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9013\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9073\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10748\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10751\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10767\ : std_logic ;
  signal \GRLFPC20.N_2403\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8302\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8356\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8675\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8242\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7965\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7905\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7729\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8293\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8332\ : std_logic ;
  signal \GRLFPC20.N_2402\ : std_logic ;
  signal \GRLFPC20.N_2074\ : std_logic ;
  signal \GRLFPC20.V.FSR.CEXC_2_SQMUXA\ : std_logic ;
  signal \GRLFPC20.V.FSR.CEXC_3_SQMUXA\ : std_logic ;
  signal \GRLFPC20.N_1837\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8788\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2693\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10724\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10154\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10166\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10170\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1101\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12021_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2818\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9828\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2335\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_967\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_969\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1580\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_972\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_991_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1006\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1006_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_830\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1009\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_796\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1011_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1012\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1267\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1034\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1347\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9946_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1187\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1014\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1036\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1041\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1047\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_838_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_841_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_836_I\ : std_logic ;
  signal \GRLFPC20.N_2361\ : std_logic ;
  signal \GRLFPC20.N_2386\ : std_logic ;
  signal \GRLFPC20.COMB.UN1_R.I.V\ : std_logic ;
  signal \GRLFPC20.N_1536\ : std_logic ;
  signal \GRLFPC20.N_1537\ : std_logic ;
  signal \GRLFPC20.N_1538\ : std_logic ;
  signal \GRLFPC20.N_2146\ : std_logic ;
  signal \GRLFPC20.N_1310\ : std_logic ;
  signal \GRLFPC20.N_1309\ : std_logic ;
  signal \GRLFPC20.N_1306\ : std_logic ;
  signal \GRLFPC20.N_1307\ : std_logic ;
  signal \GRLFPC20.N_2345\ : std_logic ;
  signal \GRLFPC20.N_2347\ : std_logic ;
  signal \GRLFPC20.N_2354\ : std_logic ;
  signal \GRLFPC20.N_2374\ : std_logic ;
  signal \GRLFPC20.N_2375\ : std_logic ;
  signal \GRLFPC20.N_2376\ : std_logic ;
  signal \GRLFPC20.N_2377\ : std_logic ;
  signal \GRLFPC20.N_2379\ : std_logic ;
  signal \GRLFPC20.N_2381\ : std_logic ;
  signal \GRLFPC20.N_2382\ : std_logic ;
  signal \GRLFPC20.N_2383\ : std_logic ;
  signal \GRLFPC20.N_2396\ : std_logic ;
  signal \GRLFPC20.N_2398\ : std_logic ;
  signal \GRLFPC20.N_2399\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_767_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_983\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_999_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1002_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1048_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1186\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1231\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2336\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_866\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1775\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12196_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_803_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2380\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_846_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1175\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_428\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_595\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_411\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_398\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_211\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_254\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2125\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_205\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_16\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2706\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2697\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1342\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2707\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9408_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2214\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2797\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2708\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_314_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9601_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7868\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7872\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.UN111_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.UN213_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.UN531_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.UN528_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.UN462_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.UN459_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.UN252_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.UN18_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.UN537_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.UN393_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.UN390_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.UN255_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.UN534_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.UN549_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.UN546_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.UN543_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.UN555_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.UN552_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.UN633_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.UN36_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN26_XZYBUSLSBS\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8313\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8314\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8316\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8318\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8216\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8691\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7689\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7691\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7692\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7693\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7694\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7696\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7697\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7698\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7702\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8709\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7704\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7705\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8712\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8713\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7709\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7711\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7713\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7714\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7716\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7718\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7720\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7721\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7723\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7725\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7726\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7727\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7732\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7733\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7734\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7738\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7865\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7867\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7869\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7870\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7873\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7874\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7875\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7878\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7879\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7880\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7881\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7882\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7883\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7885\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7887\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7889\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7890\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7892\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7893\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7896\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7899\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7901\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7902\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7903\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7908\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7909\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7910\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7914\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7925\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7927\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7928\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7929\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7930\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7933\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7934\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7938\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7940\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7941\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7945\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7947\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7949\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7950\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7952\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7953\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7954\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7956\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7959\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7961\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7962\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7963\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7968\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7969\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7970\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7974\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7717\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8273\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8275\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8278\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8279\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8281\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8282\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8286\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8287\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8288\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8289\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8290\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8294\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8295\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8300\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8304\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8308\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8319\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8322\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8325\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8326\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8327\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8334\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8351\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8354\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8360\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8631\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8635\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8637\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8639\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8640\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8642\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8643\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8644\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8645\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8648\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8650\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8651\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8655\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8657\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8659\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8660\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8664\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8666\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8667\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8668\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8669\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8671\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8672\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8673\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8678\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8679\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8680\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8638\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8662\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8684\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9066\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9068\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9071\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9072\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9074\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9076\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9080\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9081\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9082\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9085\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9089\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9092\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9095\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9096\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9097\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9100\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9106\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9108\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9112\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9119\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9121\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9126\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9128\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9132\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9134\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9136\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9140\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9141\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9142\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9145\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9149\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9152\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9155\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9156\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9157\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9160\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9166\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9168\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9172\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9179\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9181\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8972\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2823\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10790\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1561\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9445\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9435\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9548\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9661\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9629\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9846\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9840\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9941\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9896\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9957\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10290\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10284\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10405\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10332\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10479\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10647\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10576\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10648\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9642\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10839\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10948\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10082\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10090\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10678\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10699\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10690\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10449\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10446\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10460\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10309\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10305\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10304\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10292\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10299\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10300\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9922\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9928\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9855\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9860\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9652\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9655\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9660\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9511\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9496\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9497\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9494\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9495\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10819\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10824\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10827\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10834\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9558\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9549\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9454\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9451\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9453\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10605\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10619\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10616\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9964\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9968\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9974\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9664_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9576_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9915_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10752_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9788_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10860\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9739_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10087_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10293_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10759_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10765_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10746_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10694_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10696_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10671_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10670_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10624_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10629_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10631_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10584_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9723_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10592_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9906_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10437_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10383_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10343_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10236_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10243_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10246_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9919_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9916_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9855_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9726\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9669_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9637_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9560_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9509_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2129\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2219\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2224\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2772\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2645\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10130\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2502\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1593\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2343\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2208\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2559\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2563\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2565\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8110\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9428\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9473\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9596\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9709\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9801\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10225\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10237\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10448\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10458\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10457\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10442\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10365\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10310\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10294\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9782\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9786\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9799\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9779\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9794\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9785\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10535\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10155\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10156\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9716\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9720\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9719\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9409\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9385\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10609\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9969\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9604\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9605\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9601\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2161\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2167\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2341\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2162_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2337_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2377\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2379\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1748\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2734\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10441_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10297\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10161_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9887_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9366_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9800_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1726\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2512\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2235\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2210\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2220\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.UN639_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.UN636_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.UN198_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.UN195_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.UN180_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.UN138_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.UN66_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN4_NOTBINFNAN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.REEXCOVUV.UN25_LOCOV\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.REEXCOVUV.UN18_LOCOV\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8315\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8317\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8320\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8329\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8331\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8352\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8353\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8224\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7686\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7687\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7688\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7699\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7701\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7710\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7715\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7719\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7722\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7724\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7728\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7730\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7731\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7735\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7736\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7737\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7863\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7864\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7877\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7886\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7891\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7895\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7897\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7898\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7900\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7904\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7906\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7907\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7911\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7912\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7913\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7922\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7923\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7924\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7932\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7935\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7937\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7946\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7951\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7955\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7957\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7958\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7960\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7964\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7966\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7967\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7971\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7972\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7973\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8111\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8115\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8269\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8280\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8310\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8372\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8552\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8553\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8554\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8572\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8582\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8587\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8632\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8633\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8634\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8647\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8656\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8661\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8663\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8665\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8670\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8674\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8676\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8677\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8681\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8682\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8683\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8781\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8782\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8786\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8787\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8837\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9005\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9031\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9064\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9075\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9077\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9078\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9083\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9086\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9087\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9088\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9090\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9091\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9093\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9102\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9104\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9110\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9111\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9113\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9114\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9115\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9117\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9118\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9120\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9122\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9123\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9124\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9125\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9135\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9137\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9138\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9143\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9146\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9147\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9148\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9150\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9153\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9162\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9164\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9170\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9171\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9173\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9174\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9175\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9177\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9178\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9180\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9182\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9183\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9185\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12248\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9967\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12180\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10522\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12238\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10524\ : std_logic ;
  signal N_3584 : std_logic ;
  signal N_3710 : std_logic ;
  signal N_3765 : std_logic ;
  signal N_3766 : std_logic ;
  signal N_3767 : std_logic ;
  signal N_3768 : std_logic ;
  signal N_3769 : std_logic ;
  signal N_3770 : std_logic ;
  signal N_3786 : std_logic ;
  signal N_3788 : std_logic ;
  signal N_3811 : std_logic ;
  signal N_3812 : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_11\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_11\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_12\ : std_logic ;
  signal N_3825 : std_logic ;
  signal N_3826 : std_logic ;
  signal N_3827 : std_logic ;
  signal N_3880 : std_logic ;
  signal N_3881 : std_logic ;
  signal N_3882 : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_11\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_11\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_12\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_12\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_13\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_13\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_14\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_14\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_15\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_15\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_16\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_16\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_17\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_17\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_18\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_18\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_19\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_19\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_20\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_20\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_21\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_21\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_22\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_22\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_23\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_23\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_24\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_24\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_25\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_25\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_26\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_26\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_27\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_27\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_28\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_28\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_29\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_29\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_30\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_30\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_31\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_31\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_32\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_32\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_33\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_33\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_34\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_34\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_35\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_35\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_36\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_36\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_37\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_37\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_38\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_38\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_39\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_39\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_40\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_40\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_41\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_41\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_42\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_42\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_43\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_43\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_44\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_44\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_45\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_45\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_46\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_46\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_47\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_47\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_48\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_48\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_49\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_49\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_50\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_50\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_51\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_51\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_52\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_52\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_53\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_53\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_54\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_54\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_55\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_55\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_56\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_56\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_57\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6.Z_AXB2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4.Z_AXB1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21.Z_AXB2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_AXB2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18.Z_AXB1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_AXB1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_AXB2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_AXB1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_AXB2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12.Z_AXB1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8.Z_AXB2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7.Z_AXB2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36.Z_AXB2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_AXB1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33.Z_AXB2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_AXB1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_AXB2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_AXB0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_AXB1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_AXB2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27.Z_AXB2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26.Z_AXB1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26.Z_AXB2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_AXB0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_AC0_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_AC0_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_AXB1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_AC0_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_AC0_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45.Z_AXB1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44.Z_AXB2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43.Z_AXB1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_AXB2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41.Z_AXB2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39.Z_AC0_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39.Z_AC0_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_AXB1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51.Z_AC0_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51.Z_AC0_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49.Z_AXB2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48.Z_AXB0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47.Z_AXB2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_AXB1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_AXB2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_943_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54.Z_C3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53.Z_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53.Z_AXB1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53.Z_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_11\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_11\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_12\ : std_logic ;
  signal N_4325 : std_logic ;
  signal N_4327 : std_logic ;
  signal N_4328 : std_logic ;
  signal N_4331 : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL_C4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_AXB0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2963_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2966_I\ : std_logic ;
  signal N_3105_TZ : std_logic ;
  signal N_3154_TZ : std_logic ;
  signal N_6674 : std_logic ;
  signal N_6675 : std_logic ;
  signal N_6682 : std_logic ;
  signal N_6683 : std_logic ;
  signal N_6690 : std_logic ;
  signal N_6691 : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\ : std_logic ;
  signal \GRLFPC20.N_1958\ : std_logic ;
  signal \GRLFPC20.N_1502_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9748\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10223_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9857_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9490_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_7_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9911_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_A2_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10943\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_6095_A2_11_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2640\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1171\ : std_logic ;
  signal RST_I : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10055_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10484_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10788_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12045_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_591_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_593_I\ : std_logic ;
  signal \GRLFPC20.N_3022_I\ : std_logic ;
  signal \GRLFPC20.N_2961_I\ : std_logic ;
  signal \GRLFPC20.N_2941_I\ : std_logic ;
  signal \GRLFPC20.N_2929_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9288_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_871_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_870_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_3_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_678_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_676_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_680_I\ : std_logic ;
  signal N_11445 : std_logic ;
  signal \GRLFPC20.COMB.UN9_CCV_2\ : std_logic ;
  signal \GRLFPC20.COMB.WREN1_11_IV_0\ : std_logic ;
  signal \GRLFPC20.N_3082\ : std_logic ;
  signal \GRLFPC20.COMB.WREN2_11_IV_0\ : std_logic ;
  signal \GRLFPC20.COMB.WREN2_11_IV_1\ : std_logic ;
  signal \GRLFPC20.COMB.SEQERR.UN3_QNE_1_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN8_NOTAINFNAN_0\ : std_logic ;
  signal \GRLFPC20.COMB.UN1_MEXC_1_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTAINFNAN_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTAINFNAN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTBINFNAN_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1157\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN3_S_SQRT_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_6095_A2_12_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_0_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_8_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_I_18_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_6081_A2_6_0\ : std_logic ;
  signal \GRLFPC20.COMB.V.A.RF1REN_1_115_I_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN12_SRTOSTICKY_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_I_I_A2_0_O2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN3_GEN_0\ : std_logic ;
  signal \GRLFPC20.COMB.V.A.AFSR_1_0\ : std_logic ;
  signal \GRLFPC20.COMB.V.A.LD_1_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN11_WQSTSETS_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN16_NOTPROP_2336_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_154_I_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_106_I_0\ : std_logic ;
  signal \GRLFPC20.V.I.V_3_SQMUXA_0\ : std_logic ;
  signal \GRLFPC20.COMB.V.I.EXEC_18_0_29_I_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.REEXCOVUV.UN13_LOCOV_0_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.REEXCOVUV.UN13_LOCOV_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN30_CONDITIONAL_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.BUSYMULXFF.UN2_TEMP_3\ : std_logic ;
  signal \GRLFPC20.COMB.V.MK.BUSY_2_1\ : std_logic ;
  signal \GRLFPC20.COMB.V.MK.RST_1_3\ : std_logic ;
  signal NN_4 : std_logic ;
  signal \GRLFPC20.R.I.V_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_0_CY\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_0_CY\ : std_logic ;
  signal N_14162 : std_logic ;
  signal N_14163 : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8537_RETI\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RET\ : std_logic ;
  signal N_14164 : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_5_N_4_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_6_N_4_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_7_N_4_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_8_N_4_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_9_N_4_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_10_N_4_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_11_N_4_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_12_N_4_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_13_N_4_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_39_U_N_3_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_39_U_N_4_3\ : std_logic ;
  signal N_14234 : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9288_I_FAST\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_3_REP1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_8_REP1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_29_REP1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_30_REP1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_1_N_4_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_1_N_6_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_9_REP1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_7_REP1\ : std_logic ;
  signal RFI2_RD1ADDR_16 : std_logic ;
  signal RFI2_RD1ADDR_17 : std_logic ;
  signal RFI2_RD1ADDR_18 : std_logic ;
  signal RFI2_RD1ADDR_19 : std_logic ;
  signal RFI2_RD2ADDR_20 : std_logic ;
  signal RFI2_RD2ADDR_21 : std_logic ;
  signal RFI2_RD2ADDR_22 : std_logic ;
  signal RFI2_RD2ADDR_23 : std_logic ;
  signal RFI2_WRADDR_24 : std_logic ;
  signal RFI2_WRADDR_25 : std_logic ;
  signal RFI2_WRADDR_26 : std_logic ;
  signal RFI2_WRADDR_27 : std_logic ;
  signal \GRLFPC20.FPI.START_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.UN38_PCTRL_NEW_I_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.UN33_PCTRL_NEW_I_0\ : std_logic ;
  signal \GRLFPC20.FPI.RST_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3I0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3I1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1I0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1I1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1I0_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1I1_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9I0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9I1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_11\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_11\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I0_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I1_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I0_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I1_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I0_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I1_2\ : std_logic ;
  signal \GRLFPC20.N_2994_I_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.U_RDN_1_5599\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_11210_I_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_587_I_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_589_I_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN2_NOTDECODEDUNIMP_0_E\ : std_logic ;
  signal \GRLFPC20.RIN.MK.LDOP_0_E\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN3_NOTRESETORUNIMP_0_E\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.UN53_SCTRL_NEW_I_0_E\ : std_logic ;
  signal \GRLFPC20.R.MK.RST2_I_E\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_2_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_541_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_548_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_559_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8314_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8313_I\ : std_logic ;
begin
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_I_1\: MUXCY_L port map (
    DI => NN_2,
    CI => NN_3,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_N_25\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_DATA_TMP\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_I_11\: MUXCY_L port map (
    DI => NN_2,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_DATA_TMP\(2),
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_N_18\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_DATA_TMP\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_I_19\: MUXCY_L port map (
    DI => NN_2,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_DATA_TMP\(1),
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_N_11\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_DATA_TMP\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_I_27\: MUXCY_L port map (
    DI => NN_2,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_DATA_TMP\(0),
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_N_4\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_DATA_TMP\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_1\: MUXCY_L port map (
    DI => NN_2,
    CI => NN_3,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_130\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_11\: MUXCY_L port map (
    DI => NN_2,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(0),
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_123\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_19\: MUXCY_L port map (
    DI => NN_2,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(1),
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_116\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_27\: MUXCY_L port map (
    DI => NN_2,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(7),
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_109\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(8));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_35\: MUXCY_L port map (
    DI => NN_2,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(2),
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_102\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_43\: MUXCY_L port map (
    DI => NN_2,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(8),
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_95\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(9));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_51\: MUXCY_L port map (
    DI => NN_2,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(3),
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_88\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_59\: MUXCY_L port map (
    DI => NN_2,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(9),
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_81\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(10));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_67\: MUXCY_L port map (
    DI => NN_2,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(17),
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_680_I\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(18));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_75\: MUXCY_L port map (
    DI => NN_2,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(4),
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_67\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_83\: MUXCY_L port map (
    DI => NN_2,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(12),
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_60\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(13));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_91\: MUXCY_L port map (
    DI => NN_2,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(5),
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_53\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_99\: MUXCY_L port map (
    DI => NN_2,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(11),
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_676_I\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(12));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_107\: MUXCY_L port map (
    DI => NN_2,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(13),
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_39\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(14));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_115\: MUXCY_L port map (
    DI => NN_2,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(6),
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_32\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_123\: MUXCY_L port map (
    DI => NN_2,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(15),
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_25\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(16));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_131\: MUXCY_L port map (
    DI => NN_2,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(14),
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_18\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(15));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_139\: MUXCY_L port map (
    DI => NN_2,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(16),
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_11\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(17));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_147\: MUXCY_L port map (
    DI => NN_2,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(10),
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_678_I\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[64]_Z5585\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(64),
    D => \GRLFPC20.FPI.RST_0\,
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[66]_Z5586\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(66),
    D => \GRLFPC20.FPI.START_0\,
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[70]_Z5587\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(70),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(68),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[71]_Z5588\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(71),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.UN38_PCTRL_NEW_I_0\,
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[72]\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(75),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12\(75),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[74]_Z5590\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(74),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_18\(74),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[76]_Z5591\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(76),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.UN33_PCTRL_NEW_I_0\,
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[78]_Z5592\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1\(7),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[79]_Z5593\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1\(6),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[80]_Z5594\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1\(5),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[81]_Z5595\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1\(4),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[82]_Z5596\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1\(3),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[83]_Z5597\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1\(2),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[84]_Z5598\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1\(1),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[85]_Z5599\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1\(0),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[0]_Z5600\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(0),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[1]_Z5601\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(1),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[2]_Z5602\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(2),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[3]_Z5603\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(3),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[4]_Z5604\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(4),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[5]_Z5605\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(5),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(5),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[6]_Z5606\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(6),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[7]_Z5607\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(7),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[8]_Z5608\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(8),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[9]_Z5609\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(9),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(9),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[10]\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(16),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[11]_Z5611\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(11),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9288_I\,
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[12]_Z5612\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(12),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(12),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[13]_Z5613\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(13),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(13),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[14]_Z5614\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(14),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(14),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[15]_Z5615\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(15),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(15),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[17]_Z5616\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(17),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[18]_Z5617\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(18),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(18),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[19]_Z5618\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(19),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[20]_Z5619\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(20),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(20),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[21]_Z5620\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(21),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(21),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[22]_Z5621\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(22),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(22),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[23]_Z5622\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(23),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(23),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[24]_Z5623\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(24),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(24),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[25]_Z5624\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(25),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[26]_Z5625\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(26),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[27]_Z5626\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(27),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(27),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[28]_Z5627\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(28),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[29]_Z5628\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRLOI\(29),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[30]_Z5629\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRLOI\(30),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[31]_Z5630\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(31),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[32]_Z5631\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(32),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[33]_Z5632\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(33),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[34]_Z5633\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRLOI\(34),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[35]_Z5634\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(35),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(35),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[36]_Z5635\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(36),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.R.MK.BUSY_Z5636\: FDR port map (
    Q => \GRLFPC20.R.MK.BUSY\,
    D => \GRLFPC20.COMB.V.MK.BUSY_2\,
    C => clk,
    R => RST_I);
\GRLFPC20.R.MK.BUSY2_Z5637\: FDR port map (
    Q => \GRLFPC20.R.MK.BUSY2\,
    D => \GRLFPC20.COMB.V.MK.BUSY2_2\,
    C => clk,
    R => RST_I);
\GRLFPC20.R.I.EXC[0]_Z5638\: FDRE port map (
    Q => \GRLFPC20.R.I.EXC\(0),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_593_I\,
    C => clk,
    R => \GRLFPC20.N_1858\,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.EXC[1]_Z5639\: FDRE port map (
    Q => \GRLFPC20.R.I.EXC\(1),
    D => \GRLFPC20.FPO.EXC\(1),
    C => clk,
    R => \GRLFPC20.N_1858\,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.EXC[2]_Z5640\: FDRE port map (
    Q => \GRLFPC20.R.I.EXC\(2),
    D => \GRLFPC20.FPO.EXC\(2),
    C => clk,
    R => \GRLFPC20.N_1858\,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.EXC[3]_Z5641\: FDRE port map (
    Q => \GRLFPC20.R.I.EXC\(3),
    D => \GRLFPC20.FPO.EXC\(3),
    C => clk,
    R => \GRLFPC20.N_1858\,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.EXC[4]_Z5642\: FDRE port map (
    Q => \GRLFPC20.R.I.EXC\(4),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_591_I\,
    C => clk,
    R => \GRLFPC20.N_1858\,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.EXC[5]_Z5643\: FDRE port map (
    Q => \GRLFPC20.R.I.EXC\(5),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(69),
    C => clk,
    R => \GRLFPC20.N_1858\,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.INST[0]_Z5644\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(0),
    D => cpi_x_inst(0),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[1]_Z5645\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(1),
    D => cpi_x_inst(1),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[2]_Z5646\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(2),
    D => cpi_x_inst(2),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[3]_Z5647\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(3),
    D => cpi_x_inst(3),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[4]_Z5648\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(4),
    D => cpi_x_inst(4),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[5]_Z5649\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(5),
    D => cpi_x_inst(5),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[6]_Z5650\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(6),
    D => cpi_x_inst(6),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[7]_Z5651\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(7),
    D => cpi_x_inst(7),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[8]_Z5652\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(8),
    D => cpi_x_inst(8),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[9]_Z5653\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(9),
    D => cpi_x_inst(9),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[10]_Z5654\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(10),
    D => cpi_x_inst(10),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[11]_Z5655\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(11),
    D => cpi_x_inst(11),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[12]_Z5656\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(12),
    D => cpi_x_inst(12),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[13]_Z5657\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(13),
    D => cpi_x_inst(13),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[14]_Z5658\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(14),
    D => cpi_x_inst(14),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[15]_Z5659\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(15),
    D => cpi_x_inst(15),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[16]_Z5660\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(16),
    D => cpi_x_inst(16),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[17]_Z5661\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(17),
    D => cpi_x_inst(17),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[18]_Z5662\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(18),
    D => cpi_x_inst(18),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[19]_Z5663\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(19),
    D => cpi_x_inst(19),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[20]_Z5664\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(20),
    D => cpi_x_inst(20),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[21]_Z5665\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(21),
    D => cpi_x_inst(21),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[22]_Z5666\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(22),
    D => cpi_x_inst(22),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[23]_Z5667\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(23),
    D => cpi_x_inst(23),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[24]_Z5668\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(24),
    D => cpi_x_inst(24),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[25]_Z5669\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(25),
    D => cpi_x_inst(25),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[26]_Z5670\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(26),
    D => cpi_x_inst(26),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[27]_Z5671\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(27),
    D => cpi_x_inst(27),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[28]_Z5672\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(28),
    D => cpi_x_inst(28),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[29]_Z5673\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(29),
    D => cpi_x_inst(29),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[30]_Z5674\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(30),
    D => cpi_x_inst(30),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.R.I.INST[31]_Z5675\: FDRE port map (
    Q => \GRLFPC20.R.I.INST\(31),
    D => cpi_x_inst(31),
    C => clk,
    R => N_3584,
    CE => N_3710);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[63]_Z5676\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(63),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(62),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[62]_Z5677\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(62),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(61),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[61]_Z5678\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(61),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10788_I\,
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[60]_Z5679\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(60),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(59),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[59]_Z5680\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(59),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(58),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[58]_Z5681\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(58),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(57),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[57]_Z5682\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(57),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10484_I\,
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[56]_Z5683\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(56),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(55),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[55]_Z5684\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(55),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(54),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[54]_Z5685\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(54),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(53),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[53]_Z5686\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(53),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(52),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[52]_Z5687\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(52),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(51),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[51]_Z5688\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(51),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(50),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[50]_Z5689\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(50),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(49),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[49]_Z5690\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(49),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(48),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[48]_Z5691\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(48),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10055_I\,
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[47]_Z5692\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(47),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(46),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[46]_Z5693\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(46),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(45),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[45]_Z5694\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(44),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[44]_Z5695\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(43),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[43]_Z5696\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(42),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[42]_Z5697\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(41),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[41]_Z5698\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(41),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(40),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[39]_Z5699\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(39),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(38),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[38]_Z5700\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(38),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(37),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_0_Z5701\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(0),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_0_CY\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_0\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_S_0\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_0\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_0_CY\,
    O => \GRLFPC20.FPO.EXP\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_1_Z5703\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(1),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_0\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_1\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_S_1\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_1\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_0\,
    O => \GRLFPC20.FPO.EXP\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_2_Z5705\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(2),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_1\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_2\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_S_2\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_2\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_1\,
    O => \GRLFPC20.FPO.EXP\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_3_Z5707\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(3),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_2\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_3\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_S_3\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_3\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_2\,
    O => \GRLFPC20.FPO.EXP\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_4_Z5709\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(4),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_3\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_4\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_4\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_S_4\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_4\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_3\,
    O => \GRLFPC20.FPO.EXP\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_5_Z5711\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(5),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_4\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_5\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_5\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_S_5\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_5\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_4\,
    O => \GRLFPC20.FPO.EXP\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_6_Z5713\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(6),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_5\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_6\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_6\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_S_6\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_6\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_5\,
    O => \GRLFPC20.FPO.EXP\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_7_Z5715\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(7),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_6\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_7\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_7\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_S_7\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_7\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_6\,
    O => \GRLFPC20.FPO.EXP\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_8_Z5717\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(8),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_7\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_8\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_8\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_S_8\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_8\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_7\,
    O => \GRLFPC20.FPO.EXP\(8));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_9_Z5719\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(9),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_8\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_9\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_9\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_S_9\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_9\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_8\,
    O => \GRLFPC20.FPO.EXP\(9));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_10_Z5721\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(10),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_9\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_10\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_10\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_S_10\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_10\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_9\,
    O => \GRLFPC20.FPO.EXP\(10));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_11_Z5723\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(11),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_10\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_11\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_11\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_S_11\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_11\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_10\,
    O => N_3811);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_S_12\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_12\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_11\,
    O => N_3812);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_0_Z5726\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(0),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_0_CY\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_0\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_0\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_0\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_0_CY\,
    O => N_3825);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_1_Z5728\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(1),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_0\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_1\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_1\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_1\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_0\,
    O => N_3826);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_2_Z5730\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(2),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_1\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_2\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_2\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_2\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_1\,
    O => N_3827);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_3_Z5732\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(3),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_2\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_3\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_3\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_3\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_2\,
    O => \GRLFPC20.FPO.FRAC\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_4_Z5734\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(4),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_3\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_4\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_4\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_4\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_4\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_3\,
    O => \GRLFPC20.FPO.FRAC\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_5_Z5736\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(5),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_4\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_5\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_5\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_5\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_5\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_4\,
    O => \GRLFPC20.FPO.FRAC\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_6_Z5738\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(6),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_5\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_6\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_6\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_6\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_6\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_5\,
    O => \GRLFPC20.FPO.FRAC\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_7_Z5740\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(7),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_6\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_7\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_7\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_7\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_7\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_6\,
    O => \GRLFPC20.FPO.FRAC\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_8_Z5742\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(8),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_7\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_8\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_8\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_8\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_8\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_7\,
    O => \GRLFPC20.FPO.FRAC\(8));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_9_Z5744\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(9),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_8\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_9\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_9\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_9\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_9\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_8\,
    O => \GRLFPC20.FPO.FRAC\(9));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_10_Z5746\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(10),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_9\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_10\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_10\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_10\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_10\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_9\,
    O => \GRLFPC20.FPO.FRAC\(10));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_11_Z5748\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(11),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_10\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_11\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_11\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_11\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_11\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_10\,
    O => \GRLFPC20.FPO.FRAC\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_12_Z5750\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(12),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_11\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_12\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_12\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_12\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_12\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_11\,
    O => \GRLFPC20.FPO.FRAC\(12));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_13_Z5752\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(13),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_12\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_13\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_13\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_13\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_13\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_12\,
    O => \GRLFPC20.FPO.FRAC\(13));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_14_Z5754\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(14),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_13\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_14\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_14\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_14\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_14\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_13\,
    O => \GRLFPC20.FPO.FRAC\(14));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_15_Z5756\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(15),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_14\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_15\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_15\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_15\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_15\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_14\,
    O => \GRLFPC20.FPO.FRAC\(15));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_16_Z5758\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(16),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_15\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_16\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_16\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_16\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_16\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_15\,
    O => \GRLFPC20.FPO.FRAC\(16));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_17_Z5760\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(17),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_16\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_17\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_17\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_17\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_17\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_16\,
    O => \GRLFPC20.FPO.FRAC\(17));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_18_Z5762\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(18),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_17\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_18\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_18\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_18\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_18\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_17\,
    O => \GRLFPC20.FPO.FRAC\(18));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_19_Z5764\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(19),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_18\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_19\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_19\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_19\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_19\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_18\,
    O => \GRLFPC20.FPO.FRAC\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_20_Z5766\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(20),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_19\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_20\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_20\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_20\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_20\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_19\,
    O => \GRLFPC20.FPO.FRAC\(20));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_21_Z5768\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(21),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_20\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_21\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_21\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_21\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_21\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_20\,
    O => \GRLFPC20.FPO.FRAC\(21));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_22_Z5770\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(22),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_21\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_22\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_22\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_22\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_22\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_21\,
    O => \GRLFPC20.FPO.FRAC\(22));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_23_Z5772\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(23),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_22\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_23\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_23\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_23\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_23\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_22\,
    O => \GRLFPC20.FPO.FRAC\(23));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_24_Z5774\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(24),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_23\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_24\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_24\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_24\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_24\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_23\,
    O => \GRLFPC20.FPO.FRAC\(24));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_25_Z5776\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(25),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_24\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_25\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_25\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_25\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_25\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_24\,
    O => \GRLFPC20.FPO.FRAC\(25));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_26_Z5778\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(26),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_25\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_26\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_26\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_26\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_26\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_25\,
    O => \GRLFPC20.FPO.FRAC\(26));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_27_Z5780\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(27),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_26\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_27\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_27\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_27\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_27\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_26\,
    O => \GRLFPC20.FPO.FRAC\(27));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_28_Z5782\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(28),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_27\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_28\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_28\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_28\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_28\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_27\,
    O => \GRLFPC20.FPO.FRAC\(28));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_29_Z5784\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(29),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_28\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_29\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_29\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_29\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_29\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_28\,
    O => \GRLFPC20.FPO.FRAC\(29));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_30_Z5786\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(30),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_29\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_30\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_30\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_30\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_30\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_29\,
    O => \GRLFPC20.FPO.FRAC\(30));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_31_Z5788\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(31),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_30\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_31\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_31\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_31\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_31\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_30\,
    O => \GRLFPC20.FPO.FRAC\(31));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_32_Z5790\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(32),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_31\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_32\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_32\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_32\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_32\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_31\,
    O => \GRLFPC20.FPO.FRAC\(32));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_33_Z5792\: MUXCY_L port map (
    DI => N_3765,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_32\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_33\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_33\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_33\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_33\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_32\,
    O => \GRLFPC20.FPO.FRAC\(33));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_34_Z5794\: MUXCY_L port map (
    DI => N_3766,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_33\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_34\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_34\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_34\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_34\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_33\,
    O => \GRLFPC20.FPO.FRAC\(34));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_35_Z5796\: MUXCY_L port map (
    DI => N_3767,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_34\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_35\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_35\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_35\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_35\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_34\,
    O => \GRLFPC20.FPO.FRAC\(35));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_36_Z5798\: MUXCY_L port map (
    DI => N_3768,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_35\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_36\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_36\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_36\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_36\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_35\,
    O => \GRLFPC20.FPO.FRAC\(36));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_37_Z5800\: MUXCY_L port map (
    DI => N_3769,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_36\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_37\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_37\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_37\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_37\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_36\,
    O => \GRLFPC20.FPO.FRAC\(37));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_38_Z5802\: MUXCY_L port map (
    DI => N_3770,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_37\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_38\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_38\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_38\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_38\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_37\,
    O => \GRLFPC20.FPO.FRAC\(38));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_39_Z5804\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(39),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_38\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_39\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_39\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_39\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_39\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_38\,
    O => \GRLFPC20.FPO.FRAC\(39));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_40_Z5806\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(40),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_39\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_40\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_40\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_40\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_40\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_39\,
    O => \GRLFPC20.FPO.FRAC\(40));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_41_Z5808\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(41),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_40\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_41\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_41\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_41\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_41\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_40\,
    O => \GRLFPC20.FPO.FRAC\(41));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_42_Z5810\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(42),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_41\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_42\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_42\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_42\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_42\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_41\,
    O => \GRLFPC20.FPO.FRAC\(42));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_43_Z5812\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(43),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_42\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_43\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_43\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_43\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_43\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_42\,
    O => \GRLFPC20.FPO.FRAC\(43));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_44_Z5814\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(44),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_43\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_44\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_44\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_44\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_44\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_43\,
    O => \GRLFPC20.FPO.FRAC\(44));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_45_Z5816\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(45),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_44\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_45\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_45\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_45\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_45\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_44\,
    O => \GRLFPC20.FPO.FRAC\(45));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_46_Z5818\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(46),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_45\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_46\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_46\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_46\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_46\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_45\,
    O => \GRLFPC20.FPO.FRAC\(46));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_47_Z5820\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(47),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_46\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_47\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_47\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_47\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_47\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_46\,
    O => \GRLFPC20.FPO.FRAC\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_48_Z5822\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(48),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_47\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_48\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_48\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_48\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_48\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_47\,
    O => \GRLFPC20.FPO.FRAC\(48));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_49_Z5824\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(49),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_48\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_49\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_49\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_49\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_49\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_48\,
    O => \GRLFPC20.FPO.FRAC\(49));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_50_Z5826\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(50),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_49\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_50\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_50\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_50\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_50\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_49\,
    O => \GRLFPC20.FPO.FRAC\(50));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_51_Z5828\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(51),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_50\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_51\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_51\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_51\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_51\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_50\,
    O => \GRLFPC20.FPO.FRAC\(51));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_52_Z5830\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(52),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_51\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_52\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_52\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_52\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_52\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_51\,
    O => \GRLFPC20.FPO.FRAC\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_53_Z5832\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(53),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_52\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_53\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_53\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_53\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_53\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_52\,
    O => \GRLFPC20.FPO.FRAC\(53));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_54_Z5834\: MUXCY_L port map (
    DI => N_3786,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_53\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_54\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_54\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_54\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_54\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_53\,
    O => \GRLFPC20.FPO.FRAC\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_55_Z5836\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_753\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_54\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_55\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_55\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_55\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_55\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_54\,
    O => N_3880);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_56_Z5838\: MUXCY_L port map (
    DI => N_3788,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_55\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_56\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_56\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_56\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_56\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_55\,
    O => N_3881);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_S_57\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_57\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_56\,
    O => N_3882);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_0_Z5841\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(257),
    CI => NN_3,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_I\(0),
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_1_Z5842\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(256),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_0\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_1\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_S_1\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_1\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_0\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_2_Z5844\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(255),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_1\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_2\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_S_2\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_2\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_1\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_3_Z5846\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(254),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_2\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_3\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_S_3\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_3\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_2\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_4_Z5848\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(253),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_3\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_4\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_4\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_S_4\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_4\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_3\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_5_Z5850\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(252),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_4\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_5\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_5\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_S_5\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_5\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_4\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_6_Z5852\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(251),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_5\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_6\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_6\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_S_6\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_6\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_5\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_7_Z5854\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(250),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_6\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_7\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_7\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_S_7\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_7\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_6\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_8_Z5856\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(249),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_7\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_8\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_8\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_S_8\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_8\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_7\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(8));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_9_Z5858\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(248),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_8\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_9\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_9\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_S_9\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_9\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_8\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(9));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_10_Z5860\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(247),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_9\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_10\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_10\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_S_10\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_10\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_9\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(10));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_11_Z5862\: MUXCY_L port map (
    DI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(246),
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_10\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_11\,
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_11\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_S_11\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_11\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_10\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_S_12\: XORCY port map (
    LI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_12\,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CRY_11\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(12));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI3SJ51[18]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(18),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_753\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNIKS0D1[55]\: LUT5 
generic map(
  INIT => X"35CACA35"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(18),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(55),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_55\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNISLDQ[62]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(53));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNITMDQ[63]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIUNDQ[64]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(51));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIVODQ[65]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(50));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI0QDQ[66]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(49));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI1RDQ[67]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(48));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI2SDQ[68]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI3TDQ[69]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(46));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIRLEQ[70]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(45));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNISMEQ[71]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(44));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNITNEQ[72]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(43));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIUOEQ[73]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(42));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIVPEQ[74]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(41));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI0REQ[75]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(40));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI1SEQ[76]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(39));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIVQFQ[83]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(32));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIV6H01[102]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(13));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI08H01[103]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(12));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI19H01[104]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI2AH01[105]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(10));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI3BH01[106]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(9));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI4CH01[107]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(8));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI5DH01[108]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI6EH01[109]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIU6I01[110]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST_RNIDNHS[17]\: LUT4 
generic map(
  INIT => X"E2C0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST_RNIEOHS[17]\: LUT4 
generic map(
  INIT => X"E2C0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_RNI4AU51[6]\: LUT5 
generic map(
  INIT => X"FFE000E0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(6),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(17),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.EXTEND.TEMP_RNILLVS[0]\: LUT5 
generic map(
  INIT => X"47B8B847"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(115),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS_2\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN17_XZXBUS\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS_RNIF68J1[9]\: LUT5 
generic map(
  INIT => X"A695596A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8554\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8539\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(9),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_9\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS_RNIE58J1[8]\: LUT5 
generic map(
  INIT => X"A659956A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8553\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(8),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8539\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_8\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS_1_0_RNIBJBB1[7]\: LUT5 
generic map(
  INIT => X"A695596A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8552\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8539\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_7\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2_LUT6_2_RNIGSRG1[7]\: LUT5 
generic map(
  INIT => X"C93936C6"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RET\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8551\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(6),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_6\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2_LUT6_2_RNI8KRG1[0]\: LUT5 
generic map(
  INIT => X"C93936C6"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RET\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8550\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(5),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_5\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_1_LUT6_2_RNIF98E1[3]\: LUT5 
generic map(
  INIT => X"A965569A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8535\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8548\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_1_LUT6_2_RNIA23B1[3]\: LUT5 
generic map(
  INIT => X"A695596A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8547\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8534\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2_LUT6_2_RNIT04F6[1]\: LUT5 
generic map(
  INIT => X"A695596A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8546\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8533\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2_LUT6_2_RNI47591[0]\: LUT5 
generic map(
  INIT => X"A695596A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8545\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8532\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[41]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7876\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7700\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7936\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(41));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[43]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7874\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7698\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7934\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(43));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[28]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7889\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7713\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7949\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(28));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[27]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7890\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7714\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7950\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(27));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[25]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7892\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7716\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7952\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(25));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[24]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7893\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7717\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7953\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(24));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[23]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7894\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7718\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7954\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(23));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[18]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7899\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7723\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7959\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(18));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[42]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7875\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7699\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7935\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(42));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[40]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7877\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7701\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7937\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(40));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[26]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7891\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7715\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7951\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(26));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[20]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7897\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7721\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7957\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(20));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[19]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7898\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7722\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7958\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[17]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7900\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7724\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7960\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(17));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[33]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7884\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7708\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7944\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(33));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[0]\: LUT6_L 
generic map(
  INIT => X"FFF2F0F20F020002"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(116),
  I1 => \GRLFPC20.FPI.LDOP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7741\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7977\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[29]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7888\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7712\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7948\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(29));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[1]\: LUT6_L 
generic map(
  INIT => X"FFF2F0F20F020002"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(117),
  I1 => \GRLFPC20.FPI.LDOP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7740\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7976\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[2]\: LUT6_L 
generic map(
  INIT => X"FFFEF0FE0F0E000E"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(118),
  I1 => \GRLFPC20.FPI.LDOP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7739\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7975\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[12]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7905\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7729\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7965\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(12));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[44]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7873\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7697\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7933\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(44));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[39]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7878\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7702\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7938\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(39));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[37]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7880\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7704\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7940\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(37));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[36]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7881\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7705\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7941\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(36));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[32]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7885\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7709\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7945\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(32));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[30]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7887\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7711\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7947\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(30));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[21]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7896\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7720\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7956\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(21));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[16]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7901\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7725\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7961\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(16));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[15]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7902\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7726\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7962\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(15));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[14]\: LUT5_L 
generic map(
  INIT => X"FE54BA10"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7903\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7963\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7727\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(14));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[9]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7908\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7732\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7968\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(9));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[8]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7909\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7733\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7969\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(8));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[7]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7910\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7734\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7970\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[3]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7914\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7738\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7974\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[45]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7872\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7696\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7932\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(45));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[31]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7886\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7710\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7946\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(31));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[22]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7895\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7719\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7955\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(22));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[13]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7904\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7728\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7964\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(13));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[11]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7906\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7730\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7966\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[10]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7907\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7731\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7967\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(10));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[6]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7911\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7735\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7971\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[5]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7912\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7736\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7972\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[4]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7913\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7737\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7973\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[46]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7871\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7695\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7931\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(46));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[49]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7868\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7692\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7928\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(49));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[48]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7869\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7693\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7929\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(48));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[47]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7870\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7694\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7930\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[51]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7866\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7690\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7926\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(51));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[52]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7865\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7689\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7925\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[50]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7867\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7691\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7927\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(50));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[53]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7864\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7688\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7924\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(53));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[57]\: LUT6_L 
generic map(
  INIT => X"9F8F90801F0F1000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I3 => N_3825,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7979\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(57),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[41]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8646\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(41),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7700\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[43]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8644\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(43),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7698\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[28]\: LUT6 
generic map(
  INIT => X"0A3A0A0ACAFACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(28),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8659\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7713\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[27]\: LUT6 
generic map(
  INIT => X"0A3A0A0ACAFACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(27),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8660\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7714\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[25]\: LUT6 
generic map(
  INIT => X"0A3A0A0ACAFACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(25),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8662\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7716\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[23]\: LUT6 
generic map(
  INIT => X"0A3A0A0ACAFACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(23),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8664\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7718\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[20]\: LUT6 
generic map(
  INIT => X"0A3A0A0ACAFACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(20),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8667\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7721\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[18]\: LUT6 
generic map(
  INIT => X"0A3A0A0ACAFACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(18),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8669\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7723\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[42]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8645\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(42),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7699\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[40]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8647\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(40),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7701\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[26]\: LUT6 
generic map(
  INIT => X"0A3A0A0ACAFACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(26),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8661\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7715\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[24]\: LUT6 
generic map(
  INIT => X"0A3A0A0ACAFACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(24),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8663\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7717\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[19]\: LUT6 
generic map(
  INIT => X"0A3A0A0ACAFACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(19),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8668\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7722\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[17]\: LUT6 
generic map(
  INIT => X"0A3A0A0ACAFACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(17),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8670\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7724\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[55]\: LUT6_L 
generic map(
  INIT => X"FFF2F0F20F020002"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(171),
  I1 => \GRLFPC20.FPI.LDOP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7686\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7922\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(55));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[54]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7863\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7687\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7923\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[33]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8654\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(33),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7708\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[0]\: LUT6 
generic map(
  INIT => X"0A0A0A3ACACACAFA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(57),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8687\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7741\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[29]\: LUT6 
generic map(
  INIT => X"0A3A0A0ACAFACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(29),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8658\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7712\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[1]\: LUT6 
generic map(
  INIT => X"0A0A0A3ACACACAFA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(1),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8686\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7740\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[2]\: LUT6 
generic map(
  INIT => X"0A0A0A3ACACACAFA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(2),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8685\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7739\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[12]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8675\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(12),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7729\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[45]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8642\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(45),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7696\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[44]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8643\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(44),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7697\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[39]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8648\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(39),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7702\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[37]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8650\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(37),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7704\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[36]\: LUT6 
generic map(
  INIT => X"0A3A0A0ACAFACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(36),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8651\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7705\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[32]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8655\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(32),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7709\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[30]\: LUT6 
generic map(
  INIT => X"0A3A0A0ACAFACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(30),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8657\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7711\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[21]\: LUT6 
generic map(
  INIT => X"0A3A0A0ACAFACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(21),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8666\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7720\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[16]\: LUT6 
generic map(
  INIT => X"0A3A0A0ACAFACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(16),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8671\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7725\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[15]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8672\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(15),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7726\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[14]\: LUT6_L 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8673\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(14),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7727\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[9]\: LUT6 
generic map(
  INIT => X"0A0ACACA0A3ACAFA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8678\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(9),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7732\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[8]\: LUT6 
generic map(
  INIT => X"0A0ACACA0A3ACAFA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8679\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(8),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7733\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[7]\: LUT6 
generic map(
  INIT => X"0A0ACACA0A3ACAFA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8680\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7734\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[3]\: LUT6 
generic map(
  INIT => X"0A0A0A3ACACACAFA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8684\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7738\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[31]\: LUT6 
generic map(
  INIT => X"0A3A0A0ACAFACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(31),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8656\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7710\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[22]\: LUT6 
generic map(
  INIT => X"0A3A0A0ACAFACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(22),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8665\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7719\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[13]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8674\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(13),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7728\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[11]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8676\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(11),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7730\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[10]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8677\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7731\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[6]\: LUT6 
generic map(
  INIT => X"0A0ACACA0A3ACAFA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8681\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(6),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7735\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[5]\: LUT6 
generic map(
  INIT => X"0A0ACACA0A3ACAFA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8682\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(5),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7736\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[4]\: LUT6 
generic map(
  INIT => X"0A0A0A3ACACACAFA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(4),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8683\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7737\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[46]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8641\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(46),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7695\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[49]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8638\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(49),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7692\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[48]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8639\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(48),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7693\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[47]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8640\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(47),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7694\);
\GRLFPC20.COMB.V.FSR.CEXC_1_IV[0]\: LUT6_L 
generic map(
  INIT => X"FFFFCCDCFFFF0050"
)
port map (
  I0 => \GRLFPC20.N_1704\,
  I1 => \GRLFPC20.R.FSR.CEXC\(0),
  I2 => \GRLFPC20.R.I.EXC\(0),
  I3 => \GRLFPC20.COMB.V.FSR.AEXC_1_SN.N_7_MUX\,
  I4 => \GRLFPC20.COMB.V.FSR.CEXC_1_IV_1\(0),
  I5 => \GRLFPC20.V.FSR.CEXC_3_SQMUXA\,
  LO => \GRLFPC20.COMB.V.FSR.CEXC_1\(0));
\GRLFPC20.COMB.V.FSR.CEXC_1_IV[3]\: LUT6_L 
generic map(
  INIT => X"FFFFCCDCFFFF0050"
)
port map (
  I0 => \GRLFPC20.N_1704\,
  I1 => \GRLFPC20.R.FSR.CEXC\(3),
  I2 => \GRLFPC20.R.I.EXC\(3),
  I3 => \GRLFPC20.COMB.V.FSR.AEXC_1_SN.N_7_MUX\,
  I4 => \GRLFPC20.COMB.V.FSR.CEXC_1_IV_1\(3),
  I5 => \GRLFPC20.V.FSR.CEXC_3_SQMUXA\,
  LO => \GRLFPC20.COMB.V.FSR.CEXC_1\(3));
\GRLFPC20.COMB.V.FSR.CEXC_1_IV[2]\: LUT6_L 
generic map(
  INIT => X"FFFFFEFCFFFFFAF0"
)
port map (
  I0 => cpi_lddata(2),
  I1 => \GRLFPC20.R.FSR.CEXC\(2),
  I2 => \GRLFPC20.COMB.V.FSR.CEXC_1_IV_0\(2),
  I3 => \GRLFPC20.V.FSR.CEXC_2_SQMUXA\,
  I4 => \GRLFPC20.R.I.EXC_M\(2),
  I5 => \GRLFPC20.V.FSR.CEXC_3_SQMUXA\,
  LO => \GRLFPC20.COMB.V.FSR.CEXC_1\(2));
\GRLFPC20.COMB.V.FSR.CEXC_1_IV[1]\: LUT6_L 
generic map(
  INIT => X"FFFFCCDCFFFF0050"
)
port map (
  I0 => \GRLFPC20.N_1704\,
  I1 => \GRLFPC20.R.FSR.CEXC\(1),
  I2 => \GRLFPC20.R.I.EXC\(1),
  I3 => \GRLFPC20.COMB.V.FSR.AEXC_1_SN.N_7_MUX\,
  I4 => \GRLFPC20.COMB.V.FSR.CEXC_1_IV_1\(1),
  I5 => \GRLFPC20.V.FSR.CEXC_3_SQMUXA\,
  LO => \GRLFPC20.COMB.V.FSR.CEXC_1\(1));
\GRLFPC20.COMB.V.FSR.CEXC_1_IV[4]\: LUT6_L 
generic map(
  INIT => X"FFFFCCDCFFFF0050"
)
port map (
  I0 => \GRLFPC20.N_1704\,
  I1 => \GRLFPC20.R.FSR.CEXC\(4),
  I2 => \GRLFPC20.R.I.EXC\(4),
  I3 => \GRLFPC20.COMB.V.FSR.AEXC_1_SN.N_7_MUX\,
  I4 => \GRLFPC20.COMB.V.FSR.CEXC_1_IV_1\(4),
  I5 => \GRLFPC20.V.FSR.CEXC_3_SQMUXA\,
  LO => \GRLFPC20.COMB.V.FSR.CEXC_1\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[51]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8636\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(51),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7690\);
\GRLFPC20.COMB.WREN1_1\: LUT6 
generic map(
  INIT => X"55FF55FC55005500"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => \GRLFPC20.COMB.WREN1_2_M\,
  I2 => \GRLFPC20.COMB.WREN1_11_IV_0\,
  I3 => \GRLFPC20.WRADDR_0_SQMUXA\,
  I4 => \GRLFPC20.WREN1_1_SQMUXA\,
  I5 => holdn,
  O => rfi1_wren);
\GRLFPC20.COMB.WREN2_1\: LUT5 
generic map(
  INIT => X"AAFCAA00"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => \GRLFPC20.COMB.WREN2_11_IV_0\,
  I2 => \GRLFPC20.COMB.WREN2_11_IV_1\,
  I3 => \GRLFPC20.WRADDR_0_SQMUXA\,
  I4 => holdn,
  O => rfi2_wren);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[52]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8635\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(52),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7689\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[50]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8637\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(50),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7691\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[53]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8634\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(53),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7688\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[59]_Z6017\: LUT6_L 
generic map(
  INIT => X"CCCCFF0050505050"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9127\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(59),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9067\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_4_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(59));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW[7]_Z6018\: LUT6_L 
generic map(
  INIT => X"C300A5000F000F00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(8),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.U_RDN_1\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(9),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_10\(10),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.TEMP\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9260\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M[7]\: LUT6_L 
generic map(
  INIT => X"FF00FE10FD20FC30"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(50),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_28_0\(75),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_10\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_11\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8815\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8830\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES[38]\: LUT6_L 
generic map(
  INIT => X"50D872FA55DD77FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(39),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(38),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(38),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8709\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES[35]\: LUT6_L 
generic map(
  INIT => X"5072D8FA5577DDFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(35),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(36),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(35),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8712\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES[34]\: LUT6_L 
generic map(
  INIT => X"5072D8FA5577DDFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(34),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(35),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(34),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8713\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[114]_Z6023\: LUT4_L 
generic map(
  INIT => X"F011"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_25\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9132\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(114));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5[57]\: LUT6 
generic map(
  INIT => X"00000ACA0000FACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(173),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(115),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I4 => \GRLFPC20.FPI.LDOP\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8690\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7979\);
\GRLFPC20.COMB.V.FSR.AEXC_1[0]_Z6025\: LUT6_L 
generic map(
  INIT => X"BBBB8888BBB8BBB8"
)
port map (
  I0 => cpi_dbg_data(5),
  I1 => \GRLFPC20.N_1704\,
  I2 => \GRLFPC20.R.I.EXC\(0),
  I3 => \GRLFPC20.R.FSR.AEXC\(0),
  I4 => \GRLFPC20.COMB.V.FSR.AEXC_1_M0\(0),
  I5 => \GRLFPC20.COMB.V.FSR.AEXC_1_SN.N_7_MUX\,
  LO => \GRLFPC20.COMB.V.FSR.AEXC_1\(0));
\GRLFPC20.COMB.V.FSR.AEXC_1[1]_Z6026\: LUT6_L 
generic map(
  INIT => X"BBBB8888BBB8BBB8"
)
port map (
  I0 => cpi_dbg_data(6),
  I1 => \GRLFPC20.N_1704\,
  I2 => \GRLFPC20.R.I.EXC\(1),
  I3 => \GRLFPC20.R.FSR.AEXC\(1),
  I4 => \GRLFPC20.COMB.V.FSR.AEXC_1_M0\(1),
  I5 => \GRLFPC20.COMB.V.FSR.AEXC_1_SN.N_7_MUX\,
  LO => \GRLFPC20.COMB.V.FSR.AEXC_1\(1));
\GRLFPC20.COMB.V.FSR.AEXC_1[2]_Z6027\: LUT6_L 
generic map(
  INIT => X"BBBB8888BBB8BBB8"
)
port map (
  I0 => cpi_dbg_data(7),
  I1 => \GRLFPC20.N_1704\,
  I2 => \GRLFPC20.R.FSR.AEXC\(2),
  I3 => \GRLFPC20.R.I.EXC\(2),
  I4 => \GRLFPC20.COMB.V.FSR.AEXC_1_M0\(2),
  I5 => \GRLFPC20.COMB.V.FSR.AEXC_1_SN.N_7_MUX\,
  LO => \GRLFPC20.COMB.V.FSR.AEXC_1\(2));
\GRLFPC20.COMB.V.FSR.AEXC_1[3]_Z6028\: LUT6_L 
generic map(
  INIT => X"BBBB8888BBB8BBB8"
)
port map (
  I0 => cpi_dbg_data(8),
  I1 => \GRLFPC20.N_1704\,
  I2 => \GRLFPC20.R.FSR.AEXC\(3),
  I3 => \GRLFPC20.R.I.EXC\(3),
  I4 => \GRLFPC20.COMB.V.FSR.AEXC_1_M0\(3),
  I5 => \GRLFPC20.COMB.V.FSR.AEXC_1_SN.N_7_MUX\,
  LO => \GRLFPC20.COMB.V.FSR.AEXC_1\(3));
\GRLFPC20.COMB.V.FSR.AEXC_1[4]_Z6029\: LUT6_L 
generic map(
  INIT => X"BBBB8888BBB8BBB8"
)
port map (
  I0 => cpi_dbg_data(9),
  I1 => \GRLFPC20.N_1704\,
  I2 => \GRLFPC20.R.I.EXC\(4),
  I3 => \GRLFPC20.R.FSR.AEXC\(4),
  I4 => \GRLFPC20.COMB.V.FSR.AEXC_1_M0\(4),
  I5 => \GRLFPC20.COMB.V.FSR.AEXC_1_SN.N_7_MUX\,
  LO => \GRLFPC20.COMB.V.FSR.AEXC_1\(4));
\GRLFPC20.COMB.V.MK.RST_1_Z6030\: LUT6_L 
generic map(
  INIT => X"00CC04CC08CC0CCC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(50),
  I1 => \GRLFPC20.COMB.V.MK.RST_1_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_28_0\(75),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.BUSYMULXFF.UN2_TEMP_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8815\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8830\,
  LO => \GRLFPC20.COMB.V.MK.RST_1\);
\GRLFPC20.COMB.V.MK.BUSY_2_Z6031\: LUT6_L 
generic map(
  INIT => X"00CC04CC08CC0CCC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(50),
  I1 => \GRLFPC20.COMB.V.MK.BUSY_2_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_28_0\(75),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.BUSYMULXFF.UN2_TEMP_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8815\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8830\,
  LO => \GRLFPC20.COMB.V.MK.BUSY_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[41]\: LUT5 
generic map(
  INIT => X"1302DFCE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_601\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8325\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(42),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8646\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M[4]\: LUT6_L 
generic map(
  INIT => X"F0F1F0E0F2F3D0C0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(50),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_28_0\(75),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_11\(4),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8815\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_10\(4),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8830\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M[5]\: LUT6_L 
generic map(
  INIT => X"FF00FE10FD20FC30"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(50),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_28_0\(75),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_10\(5),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_11\(5),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8815\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8830\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M[0]\: LUT6_L 
generic map(
  INIT => X"F0F0F1E0F2D0F3C0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(50),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_28_0\(75),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_11\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_10\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8815\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8830\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M[3]\: LUT6_L 
generic map(
  INIT => X"FF00FE10FD20FC30"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(50),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_28_0\(75),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_10\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_11\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8815\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8830\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_14[4]_Z6037\: LUT6_L 
generic map(
  INIT => X"C000A0000C000A00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(8),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.U_RDN_1\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(9),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_10\(10),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.TEMP\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9260\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_14\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[43]\: LUT6 
generic map(
  INIT => X"EAFB6273C8D94051"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8322\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_601\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8320\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8321\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8644\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[42]\: LUT5 
generic map(
  INIT => X"8C04BF37"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_601\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8321\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(42),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8645\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[60]_Z6040\: LUT6_L 
generic map(
  INIT => X"F0F0FF00EEEEEEEE"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(60),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9126\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9066\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_4_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(60));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M[1]\: LUT6_L 
generic map(
  INIT => X"FF00FE10FD20FC30"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(50),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_28_0\(75),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_10\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_11\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8815\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8830\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M[2]\: LUT6_L 
generic map(
  INIT => X"F0F0F1E0F2D0F3C0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(50),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_28_0\(75),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_11\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_10\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8815\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8830\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M[6]\: LUT6_L 
generic map(
  INIT => X"FF00FE10FD20FC30"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(50),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_28_0\(75),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_10\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_11\(6),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8815\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8830\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[55]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8632\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(55),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7686\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0[54]\: LUT6 
generic map(
  INIT => X"0A3ACAFA0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8633\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(54),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7687\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[40]\: LUT5 
generic map(
  INIT => X"4C087F3B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_601\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8325\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(40),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8647\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[26]\: LUT3_L 
generic map(
  INIT => X"1B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(26),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(27),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8661\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[95]_Z6048\: LUT5_L 
generic map(
  INIT => X"AAF0CCCC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9091\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8972\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9031\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_4_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(95));
\GRLFPC20.COMB.V.FSR.CEXC_1_IV_1[0]_Z6049\: LUT6 
generic map(
  INIT => X"EFECECECAFA0A0A0"
)
port map (
  I0 => cpi_dbg_data(0),
  I1 => cpi_lddata(0),
  I2 => \GRLFPC20.N_1704\,
  I3 => \GRLFPC20.N_1306\,
  I4 => \GRLFPC20.N_2000\,
  I5 => \GRLFPC20.V.FSR.CEXC_2_SQMUXA\,
  O => \GRLFPC20.COMB.V.FSR.CEXC_1_IV_1\(0));
\GRLFPC20.COMB.V.FSR.CEXC_1_IV_1[3]_Z6050\: LUT6 
generic map(
  INIT => X"EFECECECAFA0A0A0"
)
port map (
  I0 => cpi_dbg_data(3),
  I1 => cpi_lddata(3),
  I2 => \GRLFPC20.N_1704\,
  I3 => \GRLFPC20.N_1309\,
  I4 => \GRLFPC20.N_2000\,
  I5 => \GRLFPC20.V.FSR.CEXC_2_SQMUXA\,
  O => \GRLFPC20.COMB.V.FSR.CEXC_1_IV_1\(3));
\GRLFPC20.COMB.V.FSR.CEXC_1_IV_1[1]_Z6051\: LUT6 
generic map(
  INIT => X"EFECECECAFA0A0A0"
)
port map (
  I0 => cpi_dbg_data(1),
  I1 => cpi_lddata(1),
  I2 => \GRLFPC20.N_1704\,
  I3 => \GRLFPC20.N_1307\,
  I4 => \GRLFPC20.N_2000\,
  I5 => \GRLFPC20.V.FSR.CEXC_2_SQMUXA\,
  O => \GRLFPC20.COMB.V.FSR.CEXC_1_IV_1\(1));
\GRLFPC20.COMB.V.FSR.CEXC_1_IV_1[4]_Z6052\: LUT6 
generic map(
  INIT => X"EFECECECAFA0A0A0"
)
port map (
  I0 => cpi_dbg_data(4),
  I1 => cpi_lddata(4),
  I2 => \GRLFPC20.N_1704\,
  I3 => \GRLFPC20.N_1310\,
  I4 => \GRLFPC20.N_2000\,
  I5 => \GRLFPC20.V.FSR.CEXC_2_SQMUXA\,
  O => \GRLFPC20.COMB.V.FSR.CEXC_1_IV_1\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[0]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => N_3881,
  I4 => N_3882,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(0),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7977\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[0]\: LUT5_L 
generic map(
  INIT => X"3210FEDC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8366\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8364\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(1),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8687\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[1]\: LUT5_L 
generic map(
  INIT => X"C480F7B3"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8362\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8364\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(1),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8686\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[2]\: LUT5_L 
generic map(
  INIT => X"3120FDEC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8362\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8364\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(3),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8685\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M_RNO_0[7]\: LUT6 
generic map(
  INIT => X"CFAACFFFCFAACF00"
)
port map (
  I0 => cpi_d_inst(12),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN3_NOTRESETORUNIMP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_0_SN_N_7_MUX\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_0_SN_N_6_MUX\,
  I5 => N_4331,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_11\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[12]\: LUT6 
generic map(
  INIT => X"F7D5B391E6C4A280"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8351\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8352\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8353\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8354\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8675\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[45]\: LUT6 
generic map(
  INIT => X"F7D5B391E6C4A280"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8318\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8319\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8320\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8321\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8642\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[44]\: LUT6 
generic map(
  INIT => X"FE76DC54BA329810"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8322\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8319\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8320\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8321\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8643\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[37]\: LUT5 
generic map(
  INIT => X"3210FEDC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8329\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8327\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(38),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8650\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[36]\: LUT5_L 
generic map(
  INIT => X"C840FB73"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8329\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8327\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(36),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8651\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[32]\: LUT5 
generic map(
  INIT => X"3210FEDC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8334\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8332\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(33),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8655\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[9]\: LUT5 
generic map(
  INIT => X"C480F7B3"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8354\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8356\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(9),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8678\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[8]\: LUT5 
generic map(
  INIT => X"3120FDEC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8356\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8358\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(9),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8679\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[7]\: LUT5 
generic map(
  INIT => X"C480F7B3"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8356\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8358\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8680\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[373]\: LUT6_L 
generic map(
  INIT => X"FEE88000FFFEE880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_C2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_113\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SCLSBS_1\(1),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_19\(0),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_25_I\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[31]\: LUT5_L 
generic map(
  INIT => X"C840FB73"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8334\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8332\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(31),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8656\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[11]\: LUT5 
generic map(
  INIT => X"C480F7B3"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8352\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8354\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(11),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8676\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[10]\: LUT5 
generic map(
  INIT => X"3120FDEC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8354\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8356\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(11),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8677\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[6]\: LUT5 
generic map(
  INIT => X"3120FDEC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8358\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8360\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8681\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[5]\: LUT5 
generic map(
  INIT => X"C480F7B3"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8358\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8360\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(5),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8682\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[4]\: LUT5_L 
generic map(
  INIT => X"3120FDEC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8360\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8362\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(5),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8683\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[3]\: LUT5_L 
generic map(
  INIT => X"C480F7B3"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8360\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8362\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(3),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8684\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8[57]_Z6075\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF88F8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN16_NOTPROP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_9\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.NOTPROP_3\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.STKGEN_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN20_STKOUT\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8_1\(57),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNO[67]\: LUT6_L 
generic map(
  INIT => X"141414141414FF00"
)
port map (
  I0 => cpi_d_inst(13),
  I1 => cpi_d_inst(19),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7596\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(67),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
  I5 => \GRLFPC20.FPI.START\,
  LO => NN_4);
\GRLFPC20.R.I.V_RNO\: LUT6_L 
generic map(
  INIT => X"CCCCCCCC0000FFF4"
)
port map (
  I0 => holdn,
  I1 => \GRLFPC20.R.I.V\,
  I2 => \GRLFPC20.N_1858\,
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.COMB.ANNULRES_1\,
  I5 => \GRLFPC20.V.I.V_3_SQMUXA\,
  LO => \GRLFPC20.R.I.V_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[46]\: LUT6 
generic map(
  INIT => X"F7D5B391E6C4A280"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8317\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8318\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8319\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8320\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8641\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_13[3]_Z6079\: LUT5_L 
generic map(
  INIT => X"C0A00C0A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(8),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.U_RDN_1\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(9),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.TEMP\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9260\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_13\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[48]\: LUT6 
generic map(
  INIT => X"F7D5B391E6C4A280"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8315\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8316\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8317\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8318\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8639\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[47]\: LUT6 
generic map(
  INIT => X"F7D5B391E6C4A280"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8316\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8317\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8318\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8319\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8640\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[58]_Z6082\: LUT6_L 
generic map(
  INIT => X"CCCCFF0050505050"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9128\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(58),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9068\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_4_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(58));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[49]\: LUT6 
generic map(
  INIT => X"F7D5B391E6C4A280"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8314\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8315\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8316\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8317\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8638\);
\GRLFPC20.COMB.V.FSR.FCC_1[0]_Z6084\: LUT6_L 
generic map(
  INIT => X"B8B8BB88BB88BB88"
)
port map (
  I0 => cpi_dbg_data(10),
  I1 => \GRLFPC20.N_1704\,
  I2 => \GRLFPC20.R.I.CC\(0),
  I3 => \GRLFPC20.COMB.V.FSR.FCC_1_M0\(0),
  I4 => \GRLFPC20.N_1837\,
  I5 => \GRLFPC20.N_2074\,
  LO => \GRLFPC20.COMB.V.FSR.FCC_1\(0));
\GRLFPC20.COMB.V.FSR.FCC_1[1]_Z6085\: LUT6_L 
generic map(
  INIT => X"B8B8BB88BB88BB88"
)
port map (
  I0 => cpi_dbg_data(11),
  I1 => \GRLFPC20.N_1704\,
  I2 => \GRLFPC20.R.I.CC\(1),
  I3 => \GRLFPC20.COMB.V.FSR.FCC_1_M0\(1),
  I4 => \GRLFPC20.N_1837\,
  I5 => \GRLFPC20.N_2074\,
  LO => \GRLFPC20.COMB.V.FSR.FCC_1\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[102]_Z6086\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(10),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(102),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9144\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(102));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[92]_Z6087\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(20),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(92),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9154\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(92));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_114_2.SUM3\: LUT5_L 
generic map(
  INIT => X"EAFE80A8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2966_I\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12044\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_114\(56),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_50\(316));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[70]_Z6089\: LUT5_L 
generic map(
  INIT => X"FF00D8D8"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(70),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(70),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9176\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(70));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[77]_Z6090\: LUT5_L 
generic map(
  INIT => X"FF00D8D8"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(77),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(77),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9169\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(77));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[107]_Z6091\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(5),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(107),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9139\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(107));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_25[0]_Z6092\: LUT6 
generic map(
  INIT => X"01177FFF0001177F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_C2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_113\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SCLSBS_1\(1),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_19\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_25\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[87]_Z6093\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(25),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(87),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9159\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(87));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[83]_Z6094\: LUT5_L 
generic map(
  INIT => X"FF00D8D8"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9163\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(83));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[24]_Z6095\: LUT6 
generic map(
  INIT => X"000FF0FF0C0CACAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8287\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_1_1\(26),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(24));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[26]_Z6096\: LUT6 
generic map(
  INIT => X"000FF0FF000AC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_1_1\(26),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_1_1\(28),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(26));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[28]_Z6097\: LUT6 
generic map(
  INIT => X"00F00FFFA0A0ACAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8281\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_1_1\(28),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(28));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[79]_Z6098\: LUT5_L 
generic map(
  INIT => X"FF00D8D8"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9167\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(79));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[81]_Z6099\: LUT5_L 
generic map(
  INIT => X"FF00D8D8"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(81),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(81),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9165\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(81));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_58_2.SUM4\: LUT6 
generic map(
  INIT => X"14BE41EBBE28EB82"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2966_I\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO2_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12044\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO0_4\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(59));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[1]\: LUT6 
generic map(
  INIT => X"FBF8CBC83B380B08"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => N_3881,
  I4 => N_3880,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(1),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7976\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[2]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(54),
  I4 => N_3880,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(2),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7975\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[85]_Z6103\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(27),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9161\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(85));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[88]_Z6104\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(24),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(88),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9158\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(88));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[113]_Z6105\: LUT6_L 
generic map(
  INIT => X"F0F0FF0044444444"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(113),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9073\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9013\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_4_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(113));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[3]\: LUT6 
generic map(
  INIT => X"3B0B3808FBCBF8C8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(53),
  I4 => \GRLFPC20.FPO.FRAC\(54),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12045\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7974\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[50]\: LUT6 
generic map(
  INIT => X"FD75B931EC64A820"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8314\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8313\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8315\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8316\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8637\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[112]_Z6108\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(112),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9134\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(112));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[110]_Z6109\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(2),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(110),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9136\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(110));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[106]_Z6110\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(6),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(106),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9140\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(106));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[105]_Z6111\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(7),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(105),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9141\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(105));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[104]_Z6112\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(8),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(104),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9142\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(104));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[101]_Z6113\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(11),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(101),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9145\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(101));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[97]_Z6114\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(97),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9149\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(97));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[94]_Z6115\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(18),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(94),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9152\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(94));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[91]_Z6116\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(21),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(91),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9155\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(91));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[90]_Z6117\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(22),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(90),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9156\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(90));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[89]_Z6118\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(23),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(89),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9157\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(89));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[86]_Z6119\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(26),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(86),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9160\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(86));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[80]_Z6120\: LUT5_L 
generic map(
  INIT => X"FF00D8D8"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9166\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(80));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[78]_Z6121\: LUT5_L 
generic map(
  INIT => X"FF00D8D8"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(78),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9168\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(78));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[74]_Z6122\: LUT5_L 
generic map(
  INIT => X"FF00D8D8"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(74),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(74),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9172\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(74));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[67]_Z6123\: LUT5_L 
generic map(
  INIT => X"FF00D8D8"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(67),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(67),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9179\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(67));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[65]_Z6124\: LUT5_L 
generic map(
  INIT => X"FF00D8D8"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(65),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(65),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9181\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(65));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[20]_Z6125\: LUT6 
generic map(
  INIT => X"00F00FFFA0A0ACAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8289\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_1_1\(20),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(20));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[18]_Z6126\: LUT6 
generic map(
  INIT => X"000FF0FF0A0ACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8293\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_1_1\(20),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(18));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[244]_Z6127\: LUT6_L 
generic map(
  INIT => X"FEFFF2FF0E000200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(27),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8587\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8572\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(244));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[53]\: LUT6 
generic map(
  INIT => X"07040F0CF7F4FFFC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8313\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_S0\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(54),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8634\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[111]_Z6129\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(111),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9135\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(111));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[109]_Z6130\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(3),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(109),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9137\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(109));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[108]_Z6131\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(4),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(108),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9138\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(108));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[103]_Z6132\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(9),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(103),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9143\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(103));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[100]_Z6133\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(12),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(100),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9146\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(100));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[99]_Z6134\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(13),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(99),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9147\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(99));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[98]_Z6135\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(14),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(98),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9148\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(98));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[96]_Z6136\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(16),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(96),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9150\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(96));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[93]_Z6137\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(19),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(93),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9153\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(93));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[84]_Z6138\: LUT6_L 
generic map(
  INIT => X"FFFF00002F202F20"
)
port map (
  I0 => rfo2_data1(28),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(84),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9162\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(84));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[82]_Z6139\: LUT5_L 
generic map(
  INIT => X"FF00D8D8"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9164\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(82));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[76]_Z6140\: LUT5_L 
generic map(
  INIT => X"FF00D8D8"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(76),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(76),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9170\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(76));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[75]_Z6141\: LUT5_L 
generic map(
  INIT => X"FF00D8D8"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(75),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(75),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9171\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(75));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[73]_Z6142\: LUT5_L 
generic map(
  INIT => X"FF00D8D8"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(73),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(73),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9173\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(73));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[72]_Z6143\: LUT5_L 
generic map(
  INIT => X"FF00D8D8"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(72),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(72),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9174\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(72));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[71]_Z6144\: LUT5_L 
generic map(
  INIT => X"FF00D8D8"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(71),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(71),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9175\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(71));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[69]_Z6145\: LUT5_L 
generic map(
  INIT => X"FF00D8D8"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(69),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(69),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9177\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(69));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[68]_Z6146\: LUT5_L 
generic map(
  INIT => X"FF00D8D8"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(68),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(68),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9178\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(68));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[66]_Z6147\: LUT5_L 
generic map(
  INIT => X"FF00D8D8"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(66),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(66),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9180\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(66));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[64]_Z6148\: LUT5_L 
generic map(
  INIT => X"FF00D8D8"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(64),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(64),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9182\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(64));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[63]_Z6149\: LUT5_L 
generic map(
  INIT => X"FF00D8D8"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(63),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(63),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9183\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(63));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[62]_Z6150\: LUT5_L 
generic map(
  INIT => X"CCF0AAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9005\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9124\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9064\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_4_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(62));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[61]_Z6151\: LUT5_L 
generic map(
  INIT => X"FF00D8D8"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(61),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(61),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9185\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(61));
\GRLFPC20.COMB.RF1REN_1[2]\: LUT6 
generic map(
  INIT => X"E2EEE2EEF3FFC0CC"
)
port map (
  I0 => N_11445,
  I1 => cpi_dbg_enable,
  I2 => cpi_dbg_fsr,
  I3 => cpi_dbg_write,
  I4 => \GRLFPC20.R.A.RF1REN\(2),
  I5 => holdn,
  O => rfi1_ren2);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M_RNO[7]\: LUT3 
generic map(
  INIT => X"E2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(53),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  I2 => N_4331,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_10\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[22]_Z6154\: LUT6 
generic map(
  INIT => X"00F00FFFCACACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8287\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8289\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(22));
\GRLFPC20.COMB.RF1REN_1[1]\: LUT6 
generic map(
  INIT => X"DF8ADF8ADFDF8A8A"
)
port map (
  I0 => cpi_dbg_enable,
  I1 => cpi_dbg_fsr,
  I2 => cpi_dbg_write,
  I3 => \GRLFPC20.COMB.V.A.RF1REN_1\(1),
  I4 => \GRLFPC20.R.A.RF1REN\(1),
  I5 => holdn,
  O => rfi1_ren1);
\GRLFPC20.COMB.RF2REN_1[1]\: LUT6 
generic map(
  INIT => X"DF8ADF8ADFDF8A8A"
)
port map (
  I0 => cpi_dbg_enable,
  I1 => cpi_dbg_fsr,
  I2 => cpi_dbg_write,
  I3 => \GRLFPC20.COMB.V.A.RF2REN_1\(1),
  I4 => \GRLFPC20.R.A.RF2REN\(1),
  I5 => holdn,
  O => rfi2_ren1);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES[56]\: LUT6_L 
generic map(
  INIT => X"FF55FE54FB51FA50"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_187\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8631\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(56),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(55),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8691\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[115]_Z6158\: LUT6_L 
generic map(
  INIT => X"F0F0CCAA00000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(115),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9071\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_4_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(115));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[36]_Z6159\: LUT6 
generic map(
  INIT => X"00F00FFFACACACAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8273\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8275\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(36));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[31]_Z6160\: LUT6 
generic map(
  INIT => X"00F00FFFCACACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8278\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8280\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(31));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[30]_Z6161\: LUT6 
generic map(
  INIT => X"00F00FFFCACACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8279\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8281\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(30));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[29]_Z6162\: LUT6 
generic map(
  INIT => X"00F00FFFACACACAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8280\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8282\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(29));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[27]_Z6163\: LUT6 
generic map(
  INIT => X"00F00FFFCACACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8282\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8284\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(27));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[25]_Z6164\: LUT6 
generic map(
  INIT => X"00F00FFFCACACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8284\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8286\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(25));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[23]_Z6165\: LUT6 
generic map(
  INIT => X"00F00FFFCACACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8286\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8288\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(23));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[21]_Z6166\: LUT6 
generic map(
  INIT => X"00F00FFFCACACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8288\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8290\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(21));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[19]_Z6167\: LUT6 
generic map(
  INIT => X"00F00FFFCACACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8290\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8292\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[17]_Z6168\: LUT6 
generic map(
  INIT => X"00F00FFFACACACAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8292\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8294\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(17));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[16]_Z6169\: LUT6 
generic map(
  INIT => X"00F00FFFACACACAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8293\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8295\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(16));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[9]_Z6170\: LUT6 
generic map(
  INIT => X"00F00FFFACACACAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8300\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8302\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(9));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[7]_Z6171\: LUT6 
generic map(
  INIT => X"00F00FFFCACACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8302\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8304\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[5]_Z6172\: LUT6 
generic map(
  INIT => X"00F00FFFACACACAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8304\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8306\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[3]_Z6173\: LUT6 
generic map(
  INIT => X"00F00FFFCACACACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8306\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8308\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[1]_Z6174\: LUT6 
generic map(
  INIT => X"000FF0FFACACACAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.LIB\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8310\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8308\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(1));
\GRLFPC20.V.FSR.CEXC_3_SQMUXA_Z6175\: LUT6 
generic map(
  INIT => X"0000000000010101"
)
port map (
  I0 => \GRLFPC20.N_1704\,
  I1 => \GRLFPC20.N_1338\,
  I2 => \GRLFPC20.N_2000\,
  I3 => \GRLFPC20.N_1837\,
  I4 => \GRLFPC20.N_2074\,
  I5 => \GRLFPC20.N_2112\,
  O => \GRLFPC20.V.FSR.CEXC_3_SQMUXA\);
\GRLFPC20.V.FSR.CEXC_2_SQMUXA_Z6176\: LUT6 
generic map(
  INIT => X"0404040404040004"
)
port map (
  I0 => \GRLFPC20.N_1704\,
  I1 => \GRLFPC20.N_1338\,
  I2 => \GRLFPC20.N_2000\,
  I3 => \GRLFPC20.N_1837\,
  I4 => \GRLFPC20.COMB.V.STATE_9\(1),
  I5 => \GRLFPC20.COMB.V.STATE_9\(0),
  O => \GRLFPC20.V.FSR.CEXC_2_SQMUXA\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[33]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(23),
  I4 => \GRLFPC20.FPO.FRAC\(24),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(33),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7944\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[41]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(15),
  I4 => \GRLFPC20.FPO.FRAC\(16),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(41),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7936\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[46]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(10),
  I4 => \GRLFPC20.FPO.FRAC\(11),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(46),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7931\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[51]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(5),
  I4 => \GRLFPC20.FPO.FRAC\(6),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(51),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7926\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[29]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(27),
  I4 => \GRLFPC20.FPO.FRAC\(28),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(29),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7948\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES[57]\: LUT6_L 
generic map(
  INIT => X"FFF7FFFFCCC4CCCC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_S0\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8690\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_2.SUM5\: LUT6 
generic map(
  INIT => X"277272278EE8E88E"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_58_2.CO1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7512\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12044\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_2.CO3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(60));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[12]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(44),
  I4 => \GRLFPC20.FPO.FRAC\(45),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(12),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7965\);
\GRLFPC20.COMB.V.FSR.AEXC_1_SN.M3\: LUT6 
generic map(
  INIT => X"5030FFFFFFFFFFFF"
)
port map (
  I0 => cpi_x_inst(19),
  I1 => \GRLFPC20.R.I.INST\(19),
  I2 => \GRLFPC20.R.X.LD\,
  I3 => \GRLFPC20.COMB.UN1_R.I.V\,
  I4 => \GRLFPC20.N_2146\,
  I5 => \GRLFPC20.N_2074\,
  O => \GRLFPC20.COMB.V.FSR.AEXC_1_SN.N_7_MUX\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[52]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(4),
  I4 => \GRLFPC20.FPO.FRAC\(5),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(52),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7925\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[50]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(6),
  I4 => \GRLFPC20.FPO.FRAC\(7),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(50),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7927\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[49]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(7),
  I4 => \GRLFPC20.FPO.FRAC\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(49),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7928\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[48]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(8),
  I4 => \GRLFPC20.FPO.FRAC\(9),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(48),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7929\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[47]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(9),
  I4 => \GRLFPC20.FPO.FRAC\(10),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(47),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7930\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[44]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(12),
  I4 => \GRLFPC20.FPO.FRAC\(13),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(44),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7933\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[43]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(13),
  I4 => \GRLFPC20.FPO.FRAC\(14),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(43),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7934\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[39]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(17),
  I4 => \GRLFPC20.FPO.FRAC\(18),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(39),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7938\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[37]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(19),
  I4 => \GRLFPC20.FPO.FRAC\(20),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(37),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7940\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[36]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(20),
  I4 => \GRLFPC20.FPO.FRAC\(21),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(36),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7941\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[32]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(24),
  I4 => \GRLFPC20.FPO.FRAC\(25),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(32),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7945\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[30]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(26),
  I4 => \GRLFPC20.FPO.FRAC\(27),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(30),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7947\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[28]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(28),
  I4 => \GRLFPC20.FPO.FRAC\(29),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(28),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7949\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[27]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(29),
  I4 => \GRLFPC20.FPO.FRAC\(30),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(27),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7950\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[25]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(31),
  I4 => \GRLFPC20.FPO.FRAC\(32),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(25),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7952\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[24]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(32),
  I4 => \GRLFPC20.FPO.FRAC\(33),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(24),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7953\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[23]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(33),
  I4 => \GRLFPC20.FPO.FRAC\(34),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(23),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7954\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[21]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(35),
  I4 => \GRLFPC20.FPO.FRAC\(36),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(21),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7956\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[18]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(38),
  I4 => \GRLFPC20.FPO.FRAC\(39),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(18),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7959\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[16]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(40),
  I4 => \GRLFPC20.FPO.FRAC\(41),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(16),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7961\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[15]\: LUT6 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(41),
  I4 => \GRLFPC20.FPO.FRAC\(42),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(15),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7962\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[14]\: LUT6 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(42),
  I4 => \GRLFPC20.FPO.FRAC\(43),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(14),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7963\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[9]\: LUT6 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(47),
  I4 => \GRLFPC20.FPO.FRAC\(48),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(9),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7968\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[8]\: LUT6 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(48),
  I4 => \GRLFPC20.FPO.FRAC\(49),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(8),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7969\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[7]\: LUT6 
generic map(
  INIT => X"FB3BCB0BF838C808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(7),
  I4 => \GRLFPC20.FPO.FRAC\(49),
  I5 => \GRLFPC20.FPO.FRAC\(50),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7970\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[55]\: LUT6_L 
generic map(
  INIT => X"D9C85140FBEA7362"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I2 => N_3826,
  I3 => N_3827,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(55),
  I5 => N_3882,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7922\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[54]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => N_3827,
  I4 => \GRLFPC20.FPO.FRAC\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(54),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7923\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[53]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(3),
  I4 => \GRLFPC20.FPO.FRAC\(4),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(53),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7924\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[45]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(11),
  I4 => \GRLFPC20.FPO.FRAC\(12),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(45),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7932\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[42]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(14),
  I4 => \GRLFPC20.FPO.FRAC\(15),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(42),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7935\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[40]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(16),
  I4 => \GRLFPC20.FPO.FRAC\(17),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(40),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7937\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[31]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(25),
  I4 => \GRLFPC20.FPO.FRAC\(26),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(31),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7946\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[26]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(30),
  I4 => \GRLFPC20.FPO.FRAC\(31),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(26),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7951\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[22]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(34),
  I4 => \GRLFPC20.FPO.FRAC\(35),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(22),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7955\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[20]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(36),
  I4 => \GRLFPC20.FPO.FRAC\(37),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(20),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7957\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[19]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(37),
  I4 => \GRLFPC20.FPO.FRAC\(38),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(19),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7958\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[17]\: LUT6 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(39),
  I4 => \GRLFPC20.FPO.FRAC\(40),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7960\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[13]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(43),
  I4 => \GRLFPC20.FPO.FRAC\(44),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(13),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7964\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[11]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(45),
  I4 => \GRLFPC20.FPO.FRAC\(46),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(11),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7966\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[10]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(46),
  I4 => \GRLFPC20.FPO.FRAC\(47),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(10),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7967\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[6]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(50),
  I4 => \GRLFPC20.FPO.FRAC\(51),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(6),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7971\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[5]\: LUT6_L 
generic map(
  INIT => X"FBCB3B0BF8C83808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(51),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(5),
  I5 => \GRLFPC20.FPO.FRAC\(52),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7972\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4[4]\: LUT6_L 
generic map(
  INIT => X"FBCBF8C83B0B3808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPO.FRAC\(52),
  I4 => \GRLFPC20.FPO.FRAC\(53),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(4),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7973\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[102]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9084\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9144\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[92]\: LUT6 
generic map(
  INIT => X"CCCCCCCCFACC0ACC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9094\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9154\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[70]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9116\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9176\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_38_U[0]\: LUT5_L 
generic map(
  INIT => X"CFAFC0A0"
)
port map (
  I0 => rfo1_data1(31),
  I1 => rfo2_data1(31),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9249\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9252\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[77]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9109\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9169\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[107]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9079\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9139\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[87]\: LUT6 
generic map(
  INIT => X"CCCCCCCCFACC0ACC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9099\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9159\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[83]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9103\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9163\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[79]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9107\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9167\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[81]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9105\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9165\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[85]\: LUT6 
generic map(
  INIT => X"CCCCCCCCFACC0ACC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9101\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9161\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[88]\: LUT6 
generic map(
  INIT => X"CCCCCCCCFACC0ACC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9098\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9158\);
\GRLFPC20.COMB.RF2REN_1[2]\: LUT6 
generic map(
  INIT => X"DF8ADF8ADFDF8A8A"
)
port map (
  I0 => cpi_dbg_enable,
  I1 => cpi_dbg_fsr,
  I2 => cpi_dbg_write,
  I3 => \GRLFPC20.COMB.V.A.RF2REN_1\(2),
  I4 => \GRLFPC20.R.A.RF2REN\(2),
  I5 => holdn,
  O => rfi2_ren2);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[114]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFC0CAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(114),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9072\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9132\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[112]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFC0CAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9074\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9134\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[110]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFC0CAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9076\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9136\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[106]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9080\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9140\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[105]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9081\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9141\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[104]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9082\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9142\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[101]\: LUT6 
generic map(
  INIT => X"CCCCCCCCFACC0ACC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9085\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9145\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[97]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9089\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9149\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[94]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9092\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9152\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[91]\: LUT6 
generic map(
  INIT => X"CCCCCCCCFACC0ACC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9095\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9155\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[90]\: LUT6 
generic map(
  INIT => X"CCCCCCCCFACC0ACC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9096\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9156\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[89]\: LUT6 
generic map(
  INIT => X"CCCCCCCCFACC0ACC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9097\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9157\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[86]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9100\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9160\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[80]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9106\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9166\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[78]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9108\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9168\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[74]\: LUT6 
generic map(
  INIT => X"CCCCCCCCFACC0ACC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9112\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9172\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[67]\: LUT6 
generic map(
  INIT => X"CCCCCCCCFACC0ACC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9119\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9179\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[65]\: LUT6 
generic map(
  INIT => X"CCCCCCCCFACC0ACC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9121\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9181\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0[95]\: LUT4 
generic map(
  INIT => X"2F20"
)
port map (
  I0 => rfo2_data1(17),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(95),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8972\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M_RNO_0[6]\: LUT6_L 
generic map(
  INIT => X"AAAAAAAA3FC0FF00"
)
port map (
  I0 => cpi_d_inst(8),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL_C4\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_0_SN_N_6_MUX\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8115\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[55]\: LUT6 
generic map(
  INIT => X"FF550F33FFFFFFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_S0\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8632\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[54]\: LUT6 
generic map(
  INIT => X"3500FF0035FFFFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_S0\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(54),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8633\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0[62]\: LUT5 
generic map(
  INIT => X"E4FFE400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I1 => \GRLFPC20.FPI.OP1\(50),
  I2 => \GRLFPC20.FPI.OP1\(53),
  I3 => \GRLFPC20.FPI.LDOP\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(62),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9005\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[111]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFC0CAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9075\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9135\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[109]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9077\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9137\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[108]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9078\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9138\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[103]\: LUT6 
generic map(
  INIT => X"CCCCCCCCFACC0ACC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9083\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9143\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[100]\: LUT6 
generic map(
  INIT => X"CCCCCCCCFACC0ACC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9086\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9146\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[99]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9087\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9147\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[98]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9088\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9148\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[96]\: LUT6 
generic map(
  INIT => X"CCCCCCCCFACC0ACC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9090\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9150\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[93]\: LUT6 
generic map(
  INIT => X"CCCCCCCCFACC0ACC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9093\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9153\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[84]\: LUT6 
generic map(
  INIT => X"CCCCCCCCFACC0ACC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9102\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9162\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[82]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9104\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9164\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[76]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9110\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9170\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[75]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9111\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9171\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[73]\: LUT6 
generic map(
  INIT => X"CCCCCCCCFACC0ACC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9113\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9173\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[72]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9114\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9174\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[71]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9115\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9175\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[69]\: LUT6 
generic map(
  INIT => X"AAAAAAAAFCAA0CAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9117\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9177\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[68]\: LUT6 
generic map(
  INIT => X"CCCCCCCCFACC0ACC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9118\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9178\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[66]\: LUT6 
generic map(
  INIT => X"CCCCCCCCFACC0ACC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9120\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9180\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[64]\: LUT6 
generic map(
  INIT => X"CCCCCCCCFACC0ACC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9122\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9182\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[63]\: LUT6 
generic map(
  INIT => X"CCCCCCCCFACC0ACC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9123\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9183\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_3[61]\: LUT6 
generic map(
  INIT => X"CCCCCCCCFACC0ACC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9125\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9185\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_I[43]\: LUT6 
generic map(
  INIT => X"FF00CCCCF0F0AAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_601\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20[2]\: LUT6 
generic map(
  INIT => X"FFFF000005330533"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(51),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8364\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20[0]\: LUT6 
generic map(
  INIT => X"FFFF0000DD0FDD0F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(53),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8366\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20[8]\: LUT6 
generic map(
  INIT => X"00FF0F0F33335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8358\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M_RNO[4]\: LUT6 
generic map(
  INIT => X"3F3FAAAA3F3FFF00"
)
port map (
  I0 => cpi_d_inst(6),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_291_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN3_NOTRESETORUNIMP\,
  I3 => N_4328,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_0_SN_N_7_MUX\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_0_SN_N_6_MUX\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_11\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN20_STKOUT_Z6292\: LUT5 
generic map(
  INIT => X"A596B7B7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SBLSBS_1\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN16_NOTPROP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO1_0\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN18_GEN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_9\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN20_STKOUT\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20[45]\: LUT6 
generic map(
  INIT => X"00FF33330F0F5555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8321\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20[10]\: LUT6 
generic map(
  INIT => X"00FF0F0F33335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8356\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20[34]\: LUT6 
generic map(
  INIT => X"00FF0F0F33335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8332\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8_1.N_12045_I\: LUT6_L 
generic map(
  INIT => X"9669699669969669"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_58_2.CO1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7512\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12044\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_2.CO3\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12045_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20[44]\: LUT6 
generic map(
  INIT => X"00FF55550F0F3333"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8322\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20[41]\: LUT6 
generic map(
  INIT => X"00FF33330F0F5555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8325\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20[40]\: LUT6 
generic map(
  INIT => X"00FF0F0F33335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8326\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20[39]\: LUT6 
generic map(
  INIT => X"00FF33330F0F5555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8327\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20[32]\: LUT6 
generic map(
  INIT => X"00FF0F0F55553333"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8334\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20[15]\: LUT6 
generic map(
  INIT => X"333300FF0F0F5555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8351\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20[12]\: LUT6 
generic map(
  INIT => X"00FF55550F0F3333"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8354\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20[37]\: LUT6 
generic map(
  INIT => X"00FF55550F0F3333"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8329\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20[35]\: LUT6 
generic map(
  INIT => X"00FF33330F0F5555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8331\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20[14]\: LUT6 
generic map(
  INIT => X"5555333300FF0F0F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8352\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20[13]\: LUT6 
generic map(
  INIT => X"00FF0F0F33335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8353\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_RNIHM0M6\: LUT5 
generic map(
  INIT => X"EAFE80A8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2966_I\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12044\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_114\(56),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(58));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL_AXBXC7\: LUT5 
generic map(
  INIT => X"6CCCCCCC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL_C4\,
  O => N_4331);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.STKGEN_3_Z6310\: LUT6 
generic map(
  INIT => X"0000010200000201"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SBLSBS_1\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO1_0\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_943_I\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN22_NOTPROP\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SCLSBS_1\(1),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.STKGEN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8_1.SUM0_1_A2\: LUT5 
generic map(
  INIT => X"95A96A56"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2966_I\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12044\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_114\(56),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8_1[57]_Z6312\: LUT6_L 
generic map(
  INIT => X"F1F1FFF1F0F0FFF0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SBLSBS_1\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO1_0\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8_1_1\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.NOTPROP_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.STKGEN_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN22_NOTPROP\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8_1\(57));
\GRLFPC20.R.STATE_RNO[1]\: LUT6_L 
generic map(
  INIT => X"50F050F040C00000"
)
port map (
  I0 => cpi_dbg_data(28),
  I1 => cpi_exack,
  I2 => rst,
  I3 => \GRLFPC20.N_1704\,
  I4 => CPO_EXC_1,
  I5 => \GRLFPC20.COMB.V.STATE_9\(1),
  LO => \GRLFPC20.COMB.V.STATE_1_IV_I\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[117]_Z6314\: LUT6_L 
generic map(
  INIT => X"CCCCAFACCCCCA0AC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(119),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(117),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => N_3881,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(117));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[118]_Z6315\: LUT6_L 
generic map(
  INIT => X"CCCCAFACCCCCA0AC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(120),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(118),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => N_3880,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(118));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[116]_Z6316\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(116),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(118),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => N_3882,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(116));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M_RNO_0[5]\: LUT5_L 
generic map(
  INIT => X"AAAA3CF0"
)
port map (
  I0 => cpi_d_inst(5),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL_C4\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_0_SN_N_6_MUX\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8114\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIIFH73_0[47]\: LUT6 
generic map(
  INIT => X"0000000000300010"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(47),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(27),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
  I3 => \GRLFPC20.FPI.LDOP\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(12),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.NOTABORTWB\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_4\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[157]_Z6319\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(157),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(159),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(16),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(157));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[139]_Z6320\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(139),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(141),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(34),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(139));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_U\: LUT6_L 
generic map(
  INIT => X"0F0003000B000300"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(57),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(56),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[133]_Z6322\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(133),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(135),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(40),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(133));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[145]_Z6323\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(145),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(147),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(28),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(145));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[146]_Z6324\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(146),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(148),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(27),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(146));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M4\: LUT6 
generic map(
  INIT => X"00FF00FF007F00FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(5),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.FPI.LDOP\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN_0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_5_0\);
\GRLFPC20.COMB.WREN129\: LUT6 
generic map(
  INIT => X"0503000000000000"
)
port map (
  I0 => cpi_x_inst(19),
  I1 => \GRLFPC20.R.I.INST\(19),
  I2 => \GRLFPC20.R.X.LD\,
  I3 => \GRLFPC20.COMB.UN1_R.I.V\,
  I4 => \GRLFPC20.N_2146\,
  I5 => \GRLFPC20.N_2074\,
  O => \GRLFPC20.N_2112\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[247]_Z6327\: LUT6_L 
generic map(
  INIT => X"FF30FFAA003000AA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(247),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.OP1\(62),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_4_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8788\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(247));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[163]_Z6328\: LUT6_L 
generic map(
  INIT => X"AAAAAAAACFCAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(163),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(165),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.FPO.FRAC\(10),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(163));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20[48]\: LUT5 
generic map(
  INIT => X"FF330F55"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8318\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[170]_Z6330\: LUT6_L 
generic map(
  INIT => X"AAAAAAAACFCAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(170),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(172),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.FPO.FRAC\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(170));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[168]_Z6331\: LUT6_L 
generic map(
  INIT => X"AAAAAAAACFCAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(168),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(170),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.FPO.FRAC\(5),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(168));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[166]_Z6332\: LUT6_L 
generic map(
  INIT => X"AAAAAAAACFCAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(166),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(168),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.FPO.FRAC\(7),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(166));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[165]_Z6333\: LUT6_L 
generic map(
  INIT => X"AAAAAAAACFCAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(165),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(167),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.FPO.FRAC\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(165));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[164]_Z6334\: LUT6_L 
generic map(
  INIT => X"AAAAAAAACFCAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(164),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(166),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.FPO.FRAC\(9),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(164));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[162]_Z6335\: LUT6_L 
generic map(
  INIT => X"AAAAAAAACFCAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(162),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(164),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.FPO.FRAC\(11),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(162));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[161]_Z6336\: LUT6_L 
generic map(
  INIT => X"AAAAAAAACFCAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(161),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(163),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.FPO.FRAC\(12),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(161));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[160]_Z6337\: LUT6_L 
generic map(
  INIT => X"AAAAAAAACFCAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(160),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(162),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.FPO.FRAC\(13),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(160));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[159]_Z6338\: LUT6_L 
generic map(
  INIT => X"AAAAAAAACFCAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(159),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(161),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.FPO.FRAC\(14),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(159));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[158]_Z6339\: LUT6_L 
generic map(
  INIT => X"AAAAAAAACFCAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(158),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(160),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.FPO.FRAC\(15),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(158));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[156]_Z6340\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(156),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(158),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(17),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(156));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[155]_Z6341\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(155),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(157),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(18),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(155));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[154]_Z6342\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(154),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(156),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(19),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(154));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[153]_Z6343\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(153),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(155),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(20),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(153));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[152]_Z6344\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(152),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(154),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(21),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(152));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[151]_Z6345\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(151),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(153),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(22),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(151));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[150]_Z6346\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(150),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(152),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(23),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(150));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[149]_Z6347\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(149),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(151),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(24),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(149));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[148]_Z6348\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(148),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(150),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(25),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(148));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[144]_Z6349\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(144),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(146),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(29),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(144));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[137]_Z6350\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(137),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(139),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(36),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(137));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[129]_Z6351\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(129),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(131),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(44),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(129));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[126]_Z6352\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(126),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(128),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(47),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(126));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[121]_Z6353\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(121),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(123),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(52),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(121));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[249]_Z6354\: LUT6_L 
generic map(
  INIT => X"FF30FFAA003000AA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(249),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.OP1\(60),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_4_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8786\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(249));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[248]_Z6355\: LUT6_L 
generic map(
  INIT => X"FF30FFAA003000AA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(248),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.OP1\(61),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_4_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8787\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(248));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[172]_Z6356\: LUT6_L 
generic map(
  INIT => X"AAAAFECEAAAA3202"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(172),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I3 => N_3826,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_14\(172),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(172));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[171]_Z6357\: LUT6_L 
generic map(
  INIT => X"FF730040FF330000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8837\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_T_3\(0),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(171));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[169]_Z6358\: LUT6_L 
generic map(
  INIT => X"AAAAAAAACFCAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(169),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(171),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.FPO.FRAC\(4),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(169));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[167]_Z6359\: LUT6_L 
generic map(
  INIT => X"AAAAAAAACFCAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(167),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(169),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.FPO.FRAC\(6),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(167));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[147]_Z6360\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(147),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(149),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(26),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(147));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[143]_Z6361\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(143),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(145),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(30),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(143));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[142]_Z6362\: LUT6_L 
generic map(
  INIT => X"AAFEAACEAA32AA02"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(142),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I4 => \GRLFPC20.FPO.FRAC\(31),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_14\(142),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(142));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[141]_Z6363\: LUT6_L 
generic map(
  INIT => X"AAFEAACEAA32AA02"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(141),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I4 => \GRLFPC20.FPO.FRAC\(32),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_14\(141),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(141));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[140]_Z6364\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(140),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(142),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(33),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(140));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[138]_Z6365\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(138),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(140),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(35),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(138));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[136]_Z6366\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(136),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(138),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(37),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(136));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[135]_Z6367\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(135),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(137),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(38),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(135));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[134]_Z6368\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(134),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(136),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(39),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(134));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[132]_Z6369\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(132),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(134),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(41),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(132));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[131]_Z6370\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(131),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(133),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(42),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(131));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[130]_Z6371\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(130),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(132),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(43),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(130));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[128]_Z6372\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(128),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(130),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(45),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(128));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[127]_Z6373\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(127),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(129),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(46),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(127));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[125]_Z6374\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(125),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(127),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(48),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(125));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[124]_Z6375\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(124),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(126),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(49),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(124));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[123]_Z6376\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(123),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(125),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(50),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(123));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[122]_Z6377\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(122),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(124),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(51),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(122));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[120]_Z6378\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(120),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(122),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(53),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(120));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[119]_Z6379\: LUT6_L 
generic map(
  INIT => X"AAAACFCAAAAAC0CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(119),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(121),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.FPO.FRAC\(54),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(119));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12[75]_Z6380\: LUT6 
generic map(
  INIT => X"44C44444C4C44444"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_26_A0_1\(75),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_1\(75),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN30_CONDITIONAL_0\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\(7),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8830\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_10[10]_Z6381\: LUT6 
generic map(
  INIT => X"FF003030FF001212"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(20),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I4 => \GRLFPC20.FPI.LDOP\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.NOTABORTWB\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_10\(10));
\GRLFPC20.COMB.LOCK_1\: LUT5 
generic map(
  INIT => X"00000010"
)
port map (
  I0 => cpi_d_annul,
  I1 => cpi_d_trap,
  I2 => \GRLFPC20.COMB.LOCKGEN.LOCKI\,
  I3 => \GRLFPC20.R.STATE\(0),
  I4 => \GRLFPC20.R.STATE\(1),
  O => cpo_ldlock);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_1_1[28]_Z6383\: LUT5 
generic map(
  INIT => X"330F0055"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_1_1\(28));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_1_1[20]_Z6384\: LUT5 
generic map(
  INIT => X"550F0033"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_1_1\(20));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_1_1[26]_Z6385\: LUT5 
generic map(
  INIT => X"0F330055"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_1_1\(26));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[59]\: LUT4 
generic map(
  INIT => X"CCAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9067\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.NOTPROP_3_Z6387\: LUT5 
generic map(
  INIT => X"FEE9977F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_C2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_113\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SCLSBS_1\(1),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.NOTPROP_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M_RNO_0[3]\: LUT6 
generic map(
  INIT => X"AA2FAA2FFF3F000F"
)
port map (
  I0 => cpi_d_inst(11),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14\(77),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN3_NOTRESETORUNIMP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  I4 => N_4327,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_0_SN_N_6_MUX\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_11\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[173]_Z6389\: LUT6_L 
generic map(
  INIT => X"32AA323202AA0202"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(173),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I3 => \GRLFPC20.FPI.LDOP\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.NOTABORTWB\,
  I5 => N_3825,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(173));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[113]\: LUT4 
generic map(
  INIT => X"AACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9013\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW[9]_Z6391\: LUT6 
generic map(
  INIT => X"FFFCAAAAFFFCFAFA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(9),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(21),
  I3 => \GRLFPC20.R.FSR.RD\(0),
  I4 => \GRLFPC20.FPI.LDOP\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.NOTABORTWB\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(9));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[60]\: LUT4 
generic map(
  INIT => X"CCAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9066\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[58]\: LUT4 
generic map(
  INIT => X"CCAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9068\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0[244]\: LUT5_L 
generic map(
  INIT => X"FC30AAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.OP2\(52),
  I3 => \GRLFPC20.FPI.OP2\(55),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8572\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[95]\: LUT4 
generic map(
  INIT => X"AACA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9031\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[62]\: LUT4 
generic map(
  INIT => X"CCAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9064\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6.Z_C4\: LUT6 
generic map(
  INIT => X"FFFFCA00CA000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.UN534_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.UN531_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.SI_120\(49),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(63));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5.Z_C4\: LUT6 
generic map(
  INIT => X"FFFFAC00AC000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.UN528_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.UN531_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.SI_119\(50),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(62));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21.Z_C4\: LUT6 
generic map(
  INIT => X"C8FE80ECFEC8EC80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.SI_78\(35),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_AXB2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(78));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_C4\: LUT6 
generic map(
  INIT => X"BEEBEBBE28828228"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_AXB1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(74));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16.Z_C4\: LUT6 
generic map(
  INIT => X"EFFEAEEA8AA80880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_AXB1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.SI_130\(39),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(73));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14.Z_C4\: LUT6 
generic map(
  INIT => X"AF8E8E0AFAE8E8A0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_C2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.SI_71\(42),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_AXB2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(71));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_C4\: LUT6 
generic map(
  INIT => X"FFFFCA00CA000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.UN555_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.UN552_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.SI_127\(42),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(70));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12.Z_C4\: LUT6 
generic map(
  INIT => X"FFFFCA00CA000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.UN552_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.UN549_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12.Z_C3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.SI_126\(43),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(69));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11.Z_C4\: LUT6 
generic map(
  INIT => X"FFFFCA00CA000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.UN549_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.UN546_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.SI_125\(44),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(68));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10.Z_C4\: LUT6 
generic map(
  INIT => X"FFFFAC00AC000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.UN543_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.UN546_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10.Z_C3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.SI_124\(45),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(67));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9.Z_C4\: LUT6 
generic map(
  INIT => X"CDDFFEEC044CC880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.SI_8\(49),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8.Z_AXB2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(66));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7.Z_C4\: LUT6 
generic map(
  INIT => X"A880FEEAFEEAA880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7.Z_C2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.SI_64\(49),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6.Z_AXB2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(64));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36.Z_C4\: LUT6 
generic map(
  INIT => X"BEEBEBBE28828228"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_AXB1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(93));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35.Z_C4\: LUT6 
generic map(
  INIT => X"EFAEFEEA8A08A880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_AXB1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.SI_149\(20),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(92));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_C4\: LUT6 
generic map(
  INIT => X"CDDFFEEC044CC880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.SI_33\(24),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33.Z_AXB2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(91));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_C4\: LUT6 
generic map(
  INIT => X"BEEBEBBE28828228"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_AXB1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(89));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_C4\: LUT6 
generic map(
  INIT => X"A8FEFEA880EAEA80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_C2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_AXB2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.SI_87\(26),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(87));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28.Z_C4\: LUT6 
generic map(
  INIT => X"A8FE80EAFEA8EA80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.SI_85\(28),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27.Z_AXB2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(85));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27.Z_C4\: LUT6 
generic map(
  INIT => X"A880FEEAFEEAA880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.SI_84\(29),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26.Z_AXB2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(84));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22.Z_C4\: LUT6 
generic map(
  INIT => X"A880FEEAFEEAA880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22.Z_C2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.SI_79\(34),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21.Z_AXB2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(79));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43.Z_C4\: LUT6 
generic map(
  INIT => X"AF8E8E0AFAE8E8A0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_C2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.SI_100\(13),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_AXB2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(100));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_C4\: LUT6 
generic map(
  INIT => X"CEEFFDDC088CC440"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_552\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.SI_41\(16),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41.Z_AXB2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(99));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41.Z_C4\: LUT6 
generic map(
  INIT => X"FFFFCA00CA000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.UN639_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.UN636_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41.Z_C3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.SI_155\(14),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(98));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40.Z_C4\: LUT6 
generic map(
  INIT => X"FFFFAC00AC000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.UN633_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.UN636_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.SI_154\(15),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(97));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37.Z_C4\: LUT6 
generic map(
  INIT => X"CDDFFEEC044CC880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.SI_36\(21),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36.Z_AXB2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(94));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_C4\: LUT6 
generic map(
  INIT => X"EEEBBBBE88822228"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51.Z_AC0_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51.Z_AC0_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.SI_108\(5),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(109));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51.Z_C4\: LUT6 
generic map(
  INIT => X"FFFEEEEAAAA88880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51.Z_AC0_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51.Z_AC0_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.SI_108\(5),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.SI_165\(4),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(108));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48.Z_C4\: LUT6 
generic map(
  INIT => X"A8FE80EAFEA8EA80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.SI_105\(8),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47.Z_AXB2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(105));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53.Z_C4\: LUT6 
generic map(
  INIT => X"EFFEAEEA8AA80880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_AXB1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.SI_167\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(110));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_49_0_A2[258]\: LUT6_L 
generic map(
  INIT => X"C60039FF39FFC600"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO0_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_114\(56),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_49\(258));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_RNIHM0M6_0\: LUT5 
generic map(
  INIT => X"95A96A56"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2966_I\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12044\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_114\(56),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8_1.SUM0_0_0_A2\: LUT6 
generic map(
  INIT => X"6996966996696996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_58_2.CO1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7512\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12044\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_2.CO3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12045\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_2_RNIR14AJ\: LUT6 
generic map(
  INIT => X"9669699669969669"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2966_I\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO2_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12044\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO0_4\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(2));
\GRLFPC20.R.A.RF2REN_RNO[2]\: LUT4_L 
generic map(
  INIT => X"00F8"
)
port map (
  I0 => cpi_d_inst(0),
  I1 => \GRLFPC20.N_1583\,
  I2 => \GRLFPC20.COMB.RS2D_1\,
  I3 => \GRLFPC20.COMB.LOCKGEN.LOCKI\,
  LO => \GRLFPC20.N_2941_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M_RNO_0[4]\: LUT6 
generic map(
  INIT => X"FE0EF202F202F202"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(56),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  I3 => N_4328,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_10\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIIFH73[47]\: LUT6 
generic map(
  INIT => X"0000000000FC0054"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(47),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(27),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
  I3 => \GRLFPC20.FPI.LDOP\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(12),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.NOTABORTWB\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[5]\: LUT5 
generic map(
  INIT => X"0F553333"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8306\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[27]\: LUT5 
generic map(
  INIT => X"0F335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8284\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[19]\: LUT5 
generic map(
  INIT => X"55330F0F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8292\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[9]\: LUT5 
generic map(
  INIT => X"0F335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8302\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[18]\: LUT5 
generic map(
  INIT => X"550F3333"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8293\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[38]\: LUT5 
generic map(
  INIT => X"0F553333"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8273\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[36]\: LUT5 
generic map(
  INIT => X"0F553333"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8275\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[33]\: LUT5 
generic map(
  INIT => X"0F335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8278\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[32]\: LUT5 
generic map(
  INIT => X"0F335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8279\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[30]\: LUT5 
generic map(
  INIT => X"0F335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8281\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[29]\: LUT5 
generic map(
  INIT => X"0F335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8282\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[25]\: LUT5 
generic map(
  INIT => X"33550F0F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8286\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[24]\: LUT5 
generic map(
  INIT => X"33550F0F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8287\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[23]\: LUT5 
generic map(
  INIT => X"33550F0F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8288\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[22]\: LUT5 
generic map(
  INIT => X"33550F0F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8289\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[21]\: LUT5 
generic map(
  INIT => X"550F3333"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8290\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[17]\: LUT5 
generic map(
  INIT => X"55330F0F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8294\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[16]\: LUT5 
generic map(
  INIT => X"330F5555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8295\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[11]\: LUT5 
generic map(
  INIT => X"0F553333"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8300\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[7]\: LUT5 
generic map(
  INIT => X"0F335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8304\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[3]\: LUT5 
generic map(
  INIT => X"0F553333"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8308\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[42]\: LUT5 
generic map(
  INIT => X"0F335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8269\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[31]\: LUT5 
generic map(
  INIT => X"0F335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8280\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_0[1]\: LUT5 
generic map(
  INIT => X"0F335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8310\);
\GRLFPC20.R.STATE_RNO[0]\: LUT6_L 
generic map(
  INIT => X"103050F000000000"
)
port map (
  I0 => cpi_dbg_data(28),
  I1 => cpi_exack,
  I2 => rst,
  I3 => \GRLFPC20.N_1704\,
  I4 => CPO_EXC_1,
  I5 => \GRLFPC20.COMB.V.STATE_9\(0),
  LO => \GRLFPC20.COMB.V.STATE_1\(0));
\GRLFPC20.COMB.V.A.AFSR_1_Z6458\: LUT6_L 
generic map(
  INIT => X"0000000010000000"
)
port map (
  I0 => cpi_d_inst(22),
  I1 => cpi_d_inst(23),
  I2 => cpi_d_inst(30),
  I3 => cpi_d_inst(31),
  I4 => \GRLFPC20.COMB.V.A.AFSR_1_0\,
  I5 => \GRLFPC20.N_1317\,
  LO => \GRLFPC20.COMB.V.A.AFSR_1\);
\GRLFPC20.COMB.V.A.LD_1_Z6459\: LUT5_L 
generic map(
  INIT => X"00001000"
)
port map (
  I0 => cpi_d_inst(21),
  I1 => cpi_d_inst(23),
  I2 => cpi_d_inst(24),
  I3 => \GRLFPC20.COMB.V.A.LD_1_1\,
  I4 => \GRLFPC20.N_1317\,
  LO => \GRLFPC20.COMB.V.A.LD_1\);
\GRLFPC20.COMB.WREN2_11_IV_1_Z6460\: LUT6 
generic map(
  INIT => X"000000004000E000"
)
port map (
  I0 => cpi_x_inst(20),
  I1 => cpi_x_inst(25),
  I2 => \GRLFPC20.N_1475\,
  I3 => \GRLFPC20.N_1958\,
  I4 => \GRLFPC20.N_2045\,
  I5 => \GRLFPC20.R.X.SEQERR\,
  O => \GRLFPC20.COMB.WREN2_11_IV_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_1[75]_Z6461\: LUT6 
generic map(
  INIT => X"FFDFAA8AF5D5A080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(49),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(48),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(51),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(52),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8822\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8825\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_1\(75));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M_RNO[2]\: LUT6 
generic map(
  INIT => X"07FFFFFF07FF0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\(5),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.OPREXCSHFT.UN3_OPREXC\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN3_NOTRESETORUNIMP\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_0_SN_N_7_MUX\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8111\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_11\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0[171]\: LUT5 
generic map(
  INIT => X"AAAABA8A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(171),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I3 => N_3827,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8837\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_2_RNIF0K69\: LUT5 
generic map(
  INIT => X"4800FF48"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2963_I\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7512\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12044\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO0_4\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"CA0035FF35FFCA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.UN534_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.UN531_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.SI_120\(49),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"36C96C93C936936C"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.SI_78\(35),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_AXB2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(21));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"6996966996696996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_AXB1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(17));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"9AA959956556A66A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_AXB1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.SI_130\(39),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(16));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"5A6969A5A596965A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_C2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.SI_71\(42),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_AXB2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(14));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"CA0035FF35FFCA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.UN555_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.UN552_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.SI_127\(42),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(13));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"CA0035FF35FFCA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.UN552_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.UN549_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12.Z_C3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.SI_126\(43),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(12));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"CA0035FF35FFCA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.UN549_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.UN546_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.SI_125\(44),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"AC0053FF53FFAC00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.UN543_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.UN546_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10.Z_C3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.SI_124\(45),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(10));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"366CC993C993366C"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.SI_8\(49),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8.Z_AXB2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(9));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"566AA995A995566A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7.Z_C2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.SI_64\(49),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6.Z_AXB2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"6996966996696996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_AXB1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(36));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"9A59A99565A6566A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_AXB1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.SI_149\(20),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(35));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"366CC993C993366C"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.SI_33\(24),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33.Z_AXB2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(34));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"6996966996696996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_AXB1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(32));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"56A9A9566A95956A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_C2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_AXB2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.SI_87\(26),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(30));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"56A96A95A956956A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.SI_85\(28),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27.Z_AXB2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(28));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"566AA995A995566A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.SI_84\(29),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26.Z_AXB2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(27));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"566AA995A995566A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22.Z_C2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.SI_79\(34),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21.Z_AXB2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(22));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"5A6969A5A596965A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_C2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.SI_100\(13),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_AXB2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(43));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"399CC663C663399C"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_552\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.SI_41\(16),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41.Z_AXB2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(42));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"CA0035FF35FFCA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.UN639_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.UN636_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41.Z_C3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.SI_155\(14),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(41));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"AC0053FF53FFAC00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.UN633_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.UN636_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.SI_154\(15),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(40));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"366CC993C993366C"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.SI_36\(21),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36.Z_AXB2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(37));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"9996666966699996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51.Z_AC0_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51.Z_AC0_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.SI_108\(5),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"AAA999955556666A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51.Z_AC0_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51.Z_AC0_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.SI_108\(5),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.SI_165\(4),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(51));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"56A96A95A956956A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.SI_105\(8),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47.Z_AXB2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(48));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"9AA959956556A66A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_AXB1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.SI_167\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(53));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_67_RNO\: LUT6 
generic map(
  INIT => X"8070080700000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_753\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(54),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(55),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_836_I\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_680_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_99_RNO\: LUT6 
generic map(
  INIT => X"0000000087878877"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\(36),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(36),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_106_I_0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_676_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_147_RNO\: LUT6 
generic map(
  INIT => X"0000000087878877"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\(33),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(33),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_154_I_0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_678_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_9[0]_Z6496\: LUT5 
generic map(
  INIT => X"2B2B033F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7498_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SALSBS_1\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN12_GEN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN10_NOTPROP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_9\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M_RNO[0]\: LUT6 
generic map(
  INIT => X"4FFF4FFFFFFF0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\(4),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\(5),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN3_NOTRESETORUNIMP\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8109\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_0_SN_N_7_MUX\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_11\(0));
\GRLFPC20.COMB.V.FSR.FTT_1_0_IV[2]\: LUT6_L 
generic map(
  INIT => X"A2A0A28000000000"
)
port map (
  I0 => rst,
  I1 => \GRLFPC20.N_1295\,
  I2 => \GRLFPC20.R.FSR.FTT\(2),
  I3 => \GRLFPC20.R.X.SEQERR\,
  I4 => \GRLFPC20.N_1421\,
  I5 => \GRLFPC20.N_3050\,
  LO => \GRLFPC20.COMB.V.FSR.FTT_1\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M_RNO[3]\: LUT6 
generic map(
  INIT => X"FFFF2E2200002E22"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(57),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  I5 => N_4327,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_10\(3));
\GRLFPC20.COMB.V.FSR.FTT_1_0_IV[1]\: LUT6_L 
generic map(
  INIT => X"AAAAAAAAA0800000"
)
port map (
  I0 => rst,
  I1 => \GRLFPC20.N_1295\,
  I2 => \GRLFPC20.R.FSR.FTT\(1),
  I3 => \GRLFPC20.N_1421\,
  I4 => \GRLFPC20.N_3050\,
  I5 => \GRLFPC20.N_2015\,
  LO => \GRLFPC20.COMB.V.FSR.FTT_1\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M_RNO_0[1]\: LUT6 
generic map(
  INIT => X"D5FFFFFFD5FF0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\(4),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\(5),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN3_NOTRESETORUNIMP\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_0_SN_N_7_MUX\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8110\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_11\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIEBH73[47]\: LUT6 
generic map(
  INIT => X"0000000000FC0054"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(47),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
  I3 => \GRLFPC20.FPI.LDOP\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(12),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.NOTABORTWB\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_4_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN_Z6503\: LUT6 
generic map(
  INIT => X"FF00FF00FFFCFF54"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(47),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(27),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
  I3 => \GRLFPC20.FPI.LDOP\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(12),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.NOTABORTWB\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_Z6504\: LUT6 
generic map(
  INIT => X"FF00FD00FD00FD00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(47),
  I1 => \GRLFPC20.FPI.LDOP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(12),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS\,
  I5 => N_3882,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN_Z6505\: LUT6 
generic map(
  INIT => X"FF00FD00FD00FD00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(47),
  I1 => \GRLFPC20.FPI.LDOP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(12),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS\,
  I5 => N_3882,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.COMB.V.FSR.FTT_1_0_IV[0]\: LUT6_L 
generic map(
  INIT => X"AAAAAAAAAAAAA080"
)
port map (
  I0 => rst,
  I1 => \GRLFPC20.N_1295\,
  I2 => \GRLFPC20.R.FSR.FTT\(0),
  I3 => \GRLFPC20.N_1421\,
  I4 => \GRLFPC20.N_2000\,
  I5 => \GRLFPC20.N_2015\,
  LO => \GRLFPC20.COMB.V.FSR.FTT_1\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.U_RDN_1[1]_Z6507\: LUT6 
generic map(
  INIT => X"FDFCDDCCFDFCFDFC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(2),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(21),
  I3 => \GRLFPC20.R.FSR.RD\(1),
  I4 => \GRLFPC20.FPI.LDOP\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.NOTABORTWB\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.U_RDN_1\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_I_34\: LUT6 
generic map(
  INIT => X"8200140014008200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(5),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(5),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12032\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_N_4\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_I_10\: LUT6 
generic map(
  INIT => X"8124184200000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(2),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12041\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_N_25\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.BUSYMULXFF.UN2_TEMP_3_Z6510\: LUT6 
generic map(
  INIT => X"0000000000000800"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(70),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(68),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14\(77),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN2_NOTDECODEDUNIMP\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.MIFROMINST\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.BUSYMULXFF.UN2_TEMP_3\);
\GRLFPC20.COMB.V.MK.RST_1_3_Z6511\: LUT6 
generic map(
  INIT => X"0000000000000080"
)
port map (
  I0 => holdn,
  I1 => \GRLFPC20.R.MK.HOLDN2\,
  I2 => \GRLFPC20.R.MK.HOLDN1\,
  I3 => \GRLFPC20.R.MK.RST\,
  I4 => \GRLFPC20.R.MK.RST2\,
  I5 => \GRLFPC20.COMB.UN1_ANNULFPU\,
  O => \GRLFPC20.COMB.V.MK.RST_1_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_114_0_A2[56]\: LUT6 
generic map(
  INIT => X"39FFC600C60039FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2966_I\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12044\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_114\(56));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.SI_118_1.CO0\: LUT6 
generic map(
  INIT => X"EBEBBEBE41821428"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO2_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2963_I\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_2.CO2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_2.CO3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_49_0_A2_RNO[258]\: LUT5 
generic map(
  INIT => X"E080FEF8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2963_I\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12044\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO0_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6.Z_C3_Z6515\: LUT5 
generic map(
  INIT => X"FEECC880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.SI_6\(51),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6.Z_C1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.SI_63\(50),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5.Z_C3_Z6516\: LUT6 
generic map(
  INIT => X"C880FEECFEECC880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_5\(52),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4.Z_C1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4.Z_AXB1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4.Z_C3_Z6517\: LUT6 
generic map(
  INIT => X"FFF6FF60F6006000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_AXB0\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4.Z_C1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_61\(52),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19.Z_C3_Z6518\: LUT6 
generic map(
  INIT => X"CF8E8E0CFCE8E8C0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.SI_19\(38),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19.Z_C1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18.Z_AXB1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18.Z_C3_Z6519\: LUT6 
generic map(
  INIT => X"CF8E8E0CFCE8E8C0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.SI_18\(39),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18.Z_C1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_AXB1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_C3_Z6520\: LUT6 
generic map(
  INIT => X"FFFFAC00AC000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.UN390_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.UN393_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.SI_74\(39),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_C3_Z6521\: LUT3 
generic map(
  INIT => X"E8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.SI_70\(43),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8.Z_C3_Z6522\: LUT5 
generic map(
  INIT => X"FEEAA880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.SI_8\(49),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.SI_65\(48),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36.Z_C3_Z6523\: LUT5 
generic map(
  INIT => X"FEEAA880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.SI_36\(21),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.SI_93\(20),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33.Z_C3_Z6524\: LUT6 
generic map(
  INIT => X"A8FE80EAFEA8EA80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_C1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.SI_33\(24),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_AXB1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_C3_Z6525\: LUT6 
generic map(
  INIT => X"F6F9F9F660909060"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(31),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.CIN_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31.Z_C1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_AXB0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_C3_Z6526\: LUT5 
generic map(
  INIT => X"EDDE8448"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.SI_28\(29),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26.Z_C3_Z6527\: LUT5 
generic map(
  INIT => X"EDDE8448"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.SI_25\(32),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_C3_Z6528\: LUT6 
generic map(
  INIT => X"EDDEEDDEEDDE8448"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.SI_24\(33),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_AC0_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_AC0_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24.Z_C3_Z6529\: LUT6 
generic map(
  INIT => X"C8FE80ECFEC8EC80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_C1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.SI_24\(33),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_AXB1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44.Z_C3_Z6530\: LUT5 
generic map(
  INIT => X"FBBAA220"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_544\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.SI_44\(13),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.SI_101\(12),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_C3_Z6531\: LUT5 
generic map(
  INIT => X"BEEB2882"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_552\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.SI_41\(16),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41.Z_C3_Z6532\: LUT5 
generic map(
  INIT => X"FBBAA220"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_552\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.SI_41\(16),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.SI_98\(15),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40.Z_C3_Z6533\: LUT6 
generic map(
  INIT => X"FFFFAC00AC000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.UN459_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.UN462_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.SI_97\(16),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39.Z_C3_Z6534\: LUT6 
generic map(
  INIT => X"EDDEEDDEEDDE8448"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.SI_38\(19),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39.Z_AC0_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39.Z_AC0_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50.Z_C3_Z6535\: LUT6 
generic map(
  INIT => X"FF96FF6996006900"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(13),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_519\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48.Z_AXB0\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.CIN_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49.Z_C1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54.Z_C3_Z6536\: LUT6 
generic map(
  INIT => X"CF4D4D0CFCD4D4C0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_457\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.SI_54\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54.Z_C1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53.Z_AXB1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL_AXBXC4\: LUT6 
generic map(
  INIT => X"AAAAAAAA6AAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  O => N_4328);
\GRLFPC20.COMB.RDD_1.M14\: LUT4_L 
generic map(
  INIT => X"4000"
)
port map (
  I0 => cpi_d_inst(22),
  I1 => cpi_d_inst(24),
  I2 => cpi_d_inst(31),
  I3 => \GRLFPC20.COMB.RDD_1.I9_MUX\,
  LO => \GRLFPC20.COMB.RDD_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNO[11]\: LUT3_L 
generic map(
  INIT => X"01"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2502\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2_1\(11),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_7\(11),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9288_I\);
\GRLFPC20.COMB.ANNULFPU_1_IV\: LUT5 
generic map(
  INIT => X"00002700"
)
port map (
  I0 => \GRLFPC20.N_1295\,
  I1 => \GRLFPC20.R.X.FPOP\,
  I2 => \GRLFPC20.R.X.SEQERR\,
  I3 => \GRLFPC20.N_1528\,
  I4 => \GRLFPC20.N_2015\,
  O => \GRLFPC20.COMB.UN1_ANNULFPU\);
\GRLFPC20.COMB.RS1V_1_IV\: LUT6 
generic map(
  INIT => X"FEFEF0F0FEEEF000"
)
port map (
  I0 => cpi_d_cnt(0),
  I1 => cpi_d_cnt(1),
  I2 => \GRLFPC20.N_878\,
  I3 => \GRLFPC20.N_940\,
  I4 => \GRLFPC20.RS1V_0_SQMUXA\,
  I5 => \GRLFPC20.RS1V_0_SQMUXA_1\,
  O => \GRLFPC20.COMB.RS1V_1\);
\GRLFPC20.R.X.AFQ_RNIUN7K1\: LUT6 
generic map(
  INIT => X"A0A0F0B000000000"
)
port map (
  I0 => \GRLFPC20.N_1295\,
  I1 => \GRLFPC20.R.X.AFQ\,
  I2 => \GRLFPC20.R.STATE\(1),
  I3 => \GRLFPC20.R.STATE\(0),
  I4 => \GRLFPC20.R.X.SEQERR\,
  I5 => \GRLFPC20.N_3050\,
  O => \GRLFPC20.COMB.V.STATE_9\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M_RNO_0[2]\: LUT3 
generic map(
  INIT => X"B8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.RESULT\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_10\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M_RNO_2[2]\: LUT6_L 
generic map(
  INIT => X"AAAAAAAAFF003FC0"
)
port map (
  I0 => cpi_d_inst(7),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_0_SN_N_6_MUX\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8111\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN_Z6545\: LUT6 
generic map(
  INIT => X"FF00FF00FFFCFF54"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(47),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
  I3 => \GRLFPC20.FPI.LDOP\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(12),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.NOTABORTWB\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNO[57]\: LUT6_L 
generic map(
  INIT => X"0000000000000007"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_291_I\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1169\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_5\(56),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_4\(56),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_8\(56),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_7_0\(56),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10484_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN_0_Z6547\: LUT6 
generic map(
  INIT => X"FFFF0000FFFFFE00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(5),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14_2\(77),
  I4 => \GRLFPC20.FPI.LDOP\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14\(77),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0_Z6548\: LUT5 
generic map(
  INIT => X"EE00EEE0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14_2\(77),
  I3 => \GRLFPC20.FPI.LDOP\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14\(77),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_122\: LUT6 
generic map(
  INIT => X"8040201008040201"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(21),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(22),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(23),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(21),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(22),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(23),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_32\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_26\: LUT6 
generic map(
  INIT => X"8020080240100401"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(8),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(6),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(7),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(8),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_116\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_18\: LUT6 
generic map(
  INIT => X"8020080240100401"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(5),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(4),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(4),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(5),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_123\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_98\: LUT6 
generic map(
  INIT => X"8040201008040201"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(18),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(19),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(20),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(18),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(19),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(20),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_53\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_82\: LUT6 
generic map(
  INIT => X"8040201008040201"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(17),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(15),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(16),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_67\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_58\: LUT6 
generic map(
  INIT => X"8020401008020401"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(13),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(12),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(14),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(12),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(13),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(14),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_88\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_42\: LUT6 
generic map(
  INIT => X"8040201008040201"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(9),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(10),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(11),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(9),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(10),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(11),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_102\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[54]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_1\(54),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(54),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0\(54),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7\(54),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9\(54),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_12\(54),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_90\: LUT6 
generic map(
  INIT => X"8020401008020401"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(40),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(39),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(41),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(39),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(40),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(41),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_60\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_50\: LUT6 
generic map(
  INIT => X"8040201008040201"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(27),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(28),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(29),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(27),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(28),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(29),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_95\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_130\: LUT6 
generic map(
  INIT => X"8040201008040201"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(48),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(49),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(50),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(48),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(49),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(50),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_25\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_114\: LUT6 
generic map(
  INIT => X"8040201008040201"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(42),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(43),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(44),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(42),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(43),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(44),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_39\);
\GRLFPC20.COMB.LOCKGEN.UN7_DEPCHECK_RNISILP\: LUT6 
generic map(
  INIT => X"1110111011100000"
)
port map (
  I0 => cpi_d_cnt(0),
  I1 => cpi_d_cnt(1),
  I2 => \GRLFPC20.COMB.FPDECODE.ST\,
  I3 => \GRLFPC20.N_1138\,
  I4 => \GRLFPC20.N_1597\,
  I5 => \GRLFPC20.N_2103\,
  O => \GRLFPC20.COMB.LOCKGEN.LOCKI\);
\GRLFPC20.COMB.ANNULRES_1_IV\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF20FF"
)
port map (
  I0 => \GRLFPC20.N_1295\,
  I1 => \GRLFPC20.R.I.EXEC\,
  I2 => \GRLFPC20.R.X.FPOP\,
  I3 => \GRLFPC20.N_1494\,
  I4 => \GRLFPC20.N_2015\,
  I5 => \GRLFPC20.R.X.SEQERR_M\,
  O => \GRLFPC20.COMB.ANNULRES_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_138\: LUT6 
generic map(
  INIT => X"8040201008040201"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(45),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(46),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(47),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(45),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(46),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(47),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_18\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_146\: LUT6 
generic map(
  INIT => X"8040201008040201"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(51),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(52),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(53),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(51),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(52),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(53),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_11\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_66\: LUT6 
generic map(
  INIT => X"8008200240041001"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(32),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(31),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(30),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(30),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(31),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(32),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_81\);
\GRLFPC20.COMB.RDD_1.M11\: LUT6 
generic map(
  INIT => X"0008100000080000"
)
port map (
  I0 => cpi_d_inst(19),
  I1 => cpi_d_inst(20),
  I2 => cpi_d_inst(21),
  I3 => cpi_d_inst(23),
  I4 => cpi_d_inst(30),
  I5 => \GRLFPC20.N_3074\,
  O => \GRLFPC20.COMB.RDD_1.I9_MUX\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_RNID0RF2_0\: LUT6 
generic map(
  INIT => X"FF2DFFD22D00D200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(368),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(5),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO0_0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO1_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5.Z_AXBXC2\: LUT6 
generic map(
  INIT => X"366CC993C993366C"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_5\(52),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4.Z_C1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4.Z_AXB1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.SI_120\(49));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4.Z_AXBXC2\: LUT6 
generic map(
  INIT => X"F609609F09F69F60"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_AXB0\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4.Z_C1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_61\(52),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.SI_119\(50));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19.Z_AXBXC2\: LUT6 
generic map(
  INIT => X"3C6969C3C396963C"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.SI_19\(38),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19.Z_C1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18.Z_AXB1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.SI_134\(35));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18.Z_AXBXC2\: LUT6 
generic map(
  INIT => X"3C6969C3C396963C"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.SI_18\(39),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18.Z_C1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_AXB1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.SI_133\(36));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_AXBXC2\: LUT6 
generic map(
  INIT => X"9669966996696996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.SI_24\(33),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_AC0_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_AC0_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.SI_140\(29));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24.Z_AXBXC2\: LUT6 
generic map(
  INIT => X"36C96C93C936936C"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_C1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.SI_24\(33),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_AXB1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.SI_139\(30));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40.Z_AXBXC2\: LUT6 
generic map(
  INIT => X"AC0053FF53FFAC00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.UN459_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.UN462_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.SI_97\(16),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.SI_155\(14));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39.Z_AXBXC2\: LUT6 
generic map(
  INIT => X"9669966996696996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.SI_38\(19),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39.Z_AC0_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39.Z_AC0_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.SI_154\(15));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50.Z_AXBXC2\: LUT6 
generic map(
  INIT => X"9669699669969669"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(13),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_519\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48.Z_AXB0\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.CIN_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49.Z_C1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.SI_165\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48.Z_AXBXC2\: LUT3 
generic map(
  INIT => X"96"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.SI_105\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.SI_163\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55.Z_AXBXC2\: LUT5 
generic map(
  INIT => X"C663399C"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_453\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.SI_55\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.SI_112\(1),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SCLSBS_1\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54.Z_AXBXC2\: LUT6 
generic map(
  INIT => X"3C9696C3C369693C"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_457\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.SI_54\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54.Z_C1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53.Z_AXB1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL_AXBXC3\: LUT5 
generic map(
  INIT => X"CCCC6CCC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  O => N_4327);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL_AC0_5\: LUT5 
generic map(
  INIT => X"00008000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL_C4\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[48]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10154\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10157\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(48),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_1\(48),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7\(48),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(48),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(48));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.SI_118_1.SUM0\: LUT6 
generic map(
  INIT => X"6996966996696996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO2_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2963_I\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_2.CO2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.SI_118\(51));
\GRLFPC20.R.A.RF1REN_RNO_0[1]\: LUT6 
generic map(
  INIT => X"000080803320B3A0"
)
port map (
  I0 => cpi_d_inst(14),
  I1 => \GRLFPC20.N_940\,
  I2 => \GRLFPC20.N_1583\,
  I3 => \GRLFPC20.N_2512\,
  I4 => \GRLFPC20.COMB.FPDECODE.RS1D5\,
  I5 => \GRLFPC20.RS1D_CNST\,
  O => \GRLFPC20.COMB.V.A.RF1REN_1_115_I_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_3_I_Z6585\: LUT6 
generic map(
  INIT => X"0FFFC333C333A555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(174),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SS0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_3_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL[3]_Z6586\: LUT6 
generic map(
  INIT => X"ECEC2C2CECE02C20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(241),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_93\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20.V.STATE_2_SQMUXA_Z6587\: LUT6 
generic map(
  INIT => X"AAAAFFBF00000000"
)
port map (
  I0 => \GRLFPC20.N_1295\,
  I1 => \GRLFPC20.R.X.AFQ\,
  I2 => \GRLFPC20.R.STATE\(1),
  I3 => \GRLFPC20.R.STATE\(0),
  I4 => \GRLFPC20.R.X.SEQERR\,
  I5 => \GRLFPC20.N_3050\,
  O => \GRLFPC20.V.STATE_2_SQMUXA\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_18[75]\: LUT6 
generic map(
  INIT => X"EDEEEDDD21222111"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(48),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(51),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(12),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(52),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8821\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8822\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M_RNO[1]\: LUT6 
generic map(
  INIT => X"FFFFEEEC0000EEEC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.RESULT_IV_0\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS\,
  I3 => N_3812,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  I5 => N_4325,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_10\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M_RNO_1[1]\: LUT6_L 
generic map(
  INIT => X"FFFFBFAA000080AA"
)
port map (
  I0 => cpi_d_inst(9),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(63),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14_2\(77),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.TEMP_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  I5 => N_4325,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8110\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNO[48]\: LUT4_L 
generic map(
  INIT => X"0001"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2343\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_5\(47),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_7\(47),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2_1\(47),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10055_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[58]\: LUT5_L 
generic map(
  INIT => X"FFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1971\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(58),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9\(58),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7\(58),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8\(58),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(58));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[33]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFF8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9915_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9855_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2343\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7_0\(33),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(33),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9\(33),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(33));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[32]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFF2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9857_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_125\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0\(32),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(32),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(32),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8\(32),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(32));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_10\: LUT6 
generic map(
  INIT => X"8040080420100201"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(2),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN17_XZXBUS\(1),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN17_XZXBUS\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_130\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[51]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFF4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2730\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1650\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_4_1\(51),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_1\(51),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(51),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(51));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[52]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFF8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_2_0\(52),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2454_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(52),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_0\(52),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3\(52),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_11\(52),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[17]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1711\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1648\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1710\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_0\(17),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1661\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_1\(17),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(17));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_34\: LUT6 
generic map(
  INIT => X"8040201008040201"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(24),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(25),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(26),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(24),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(25),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(26),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_109\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_154_I_0_Z6600\: LUT6_L 
generic map(
  INIT => X"78787788FFFFFFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\(34),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(34),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_841_I\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_154_I_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_106_I_0_Z6601\: LUT6_L 
generic map(
  INIT => X"78787788FFFFFFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\(37),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(37),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_838_I\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_106_I_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNICSNC3[60]\: LUT6 
generic map(
  INIT => X"C3A5FFFF3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO0_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7512\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNICSNC3_0[60]\: LUT6 
generic map(
  INIT => X"3C5A000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO0_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO2_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIQNCS3[22]\: LUT6 
generic map(
  INIT => X"53FF000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SBLSBS_2\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN18_GEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6.Z_C2_Z6605\: LUT6 
generic map(
  INIT => X"FFF2FF20F2002000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(318),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(55),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.CIN_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.SI_6\(51),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21.Z_C2_Z6606\: LUT6 
generic map(
  INIT => X"FFF2FF20F2002000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(333),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(40),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.CIN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.SI_21\(36),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_C2_Z6607\: LUT6 
generic map(
  INIT => X"FF2DFFD22D00D200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(331),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(42),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.CIN_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.CIN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_C2_Z6608\: LUT6 
generic map(
  INIT => X"FF2DFFD22D00D200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(328),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(45),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.CIN_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.CIN_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_AXB2_Z6609\: LUT5 
generic map(
  INIT => X"53FFAC00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.UN390_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.UN393_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.SI_74\(39),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_AXB2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16.Z_C2_Z6610\: LUT6 
generic map(
  INIT => X"FFF2FF20F2002000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(328),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(45),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.CIN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.CIN_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.SI_16\(41),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14.Z_C2_Z6611\: LUT6 
generic map(
  INIT => X"FFF2FF20F2002000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(326),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(47),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.CIN_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.SI_14\(43),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_C2_Z6612\: LUT6 
generic map(
  INIT => X"FF2DFFD22D00D200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(324),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.CIN_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.CIN_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_AXB2_Z6613\: LUT6 
generic map(
  INIT => X"F20D20DF0DF2DF20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(324),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.CIN_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.CIN_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12.Z_AXB1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_AXB2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12.Z_C2_Z6614\: LUT6 
generic map(
  INIT => X"FFF2FF20F2002000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(324),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.CIN_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.CIN_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.SI_12\(45),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10.Z_C2_Z6615\: LUT6 
generic map(
  INIT => X"FFFFAC00AC000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.UN195_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.UN198_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10.Z_C1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.SI_10\(47),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7.Z_C2_Z6616\: LUT6 
generic map(
  INIT => X"FF2DFFD22D00D200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(318),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(55),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.CIN_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7.Z_AXB2_Z6617\: LUT4 
generic map(
  INIT => X"6996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.SI_6\(51),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7.Z_AXB2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35.Z_C2_Z6618\: LUT6 
generic map(
  INIT => X"FF2DFFD22D00D200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(346),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(27),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.CIN_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_C2_Z6619\: LUT6 
generic map(
  INIT => X"FFF2FF20F2002000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(346),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(27),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.CIN_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.SI_34\(23),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_AXB2_Z6620\: LUT5 
generic map(
  INIT => X"96696996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(31),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.CIN_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31.Z_C1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_AXB0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_AXB2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_C2_Z6621\: LUT6 
generic map(
  INIT => X"FFF2FF20F2002000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(342),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(31),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.CIN_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.CIN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.SI_30\(27),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_C2_Z6622\: LUT6 
generic map(
  INIT => X"FFFFAC00AC000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.UN252_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.UN255_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_C1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.SI_29\(28),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27.Z_C2_Z6623\: LUT6 
generic map(
  INIT => X"FF2DFFD22D00D200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(338),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(35),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.CIN_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.CIN_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27.Z_AXB2_Z6624\: LUT6 
generic map(
  INIT => X"F2200DDF0DDFF220"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(338),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(35),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.CIN_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.CIN_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26.Z_AXB1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27.Z_AXB2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26.Z_C2_Z6625\: LUT6 
generic map(
  INIT => X"FFF2FF20F2002000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(338),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(35),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.CIN_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.CIN_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.SI_26\(31),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22.Z_C2_Z6626\: LUT6 
generic map(
  INIT => X"FF2DFFD22D00D200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(333),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(40),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.CIN_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45.Z_C2_Z6627\: LUT6 
generic map(
  INIT => X"F2FF20FF00F20020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(357),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(16),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_541\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.CIN_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.SI_45\(12),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44.Z_AXB2_Z6628\: LUT6 
generic map(
  INIT => X"F2200DDF0DDFF220"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(355),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(18),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.CIN_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.CIN_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43.Z_AXB1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44.Z_AXB2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43.Z_C2_Z6629\: LUT6 
generic map(
  INIT => X"F2FF20FF00F20020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(355),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(18),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_548\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.SI_43\(14),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_C2_Z6630\: LUT6 
generic map(
  INIT => X"2DFFD2FF002D00D2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(353),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(20),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_550\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.CIN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41.Z_AXB2_Z6631\: LUT6 
generic map(
  INIT => X"E11E87781EE17887"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(21),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(21),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_554\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.CIN_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.SI_40\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41.Z_AXB2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37.Z_C2_Z6632\: LUT6 
generic map(
  INIT => X"FFF2FF20F2002000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(349),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(24),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.CIN_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.CIN_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.SI_37\(20),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_C2_Z6633\: LUT6 
generic map(
  INIT => X"2DFFD2FF002D00D2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(363),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(10),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_513\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50.Z_C2_Z6634\: LUT6 
generic map(
  INIT => X"FFFFAC00AC000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_811_I\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_812_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50.Z_C1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.SI_50\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49.Z_C2_Z6635\: LUT4 
generic map(
  INIT => X"7B12"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(13),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_519\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48.Z_AXB0\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49.Z_AXB2_Z6636\: LUT6 
generic map(
  INIT => X"E1871E781E78E187"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(13),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(13),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_521\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.CIN_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.CIN_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.SI_48\(9),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49.Z_AXB2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47.Z_C2_Z6637\: LUT6 
generic map(
  INIT => X"F2FF20FF00F20020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(359),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(14),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_523\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.CIN_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.SI_47\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_C2_Z6638\: LUT6 
generic map(
  INIT => X"2DFFD2FF002D00D2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(357),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(16),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_537\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.CIN_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_AXB2_Z6639\: LUT6 
generic map(
  INIT => X"F2200DDF0DDFF220"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(357),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(16),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.CIN_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.CIN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45.Z_AXB1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_AXB2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI3CFC3[368]\: LUT6 
generic map(
  INIT => X"FFF2FF20F2002000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(368),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(5),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.SI_56\(1),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53.Z_C2_Z6641\: LUT6 
generic map(
  INIT => X"2DFFD2FF002D00D2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(364),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(9),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_499\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[62]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFCC80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10927_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_722\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10943\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10925\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(62),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(62));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_2_Z6643\: LUT6 
generic map(
  INIT => X"F2A2C08000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1086\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8198\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8199\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8200\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8_1_1[57]_Z6644\: LUT5 
generic map(
  INIT => X"FFF2F2F2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(315),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8_0_0\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN10_NOTPROP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8_1_1\(57));
\GRLFPC20.WRDATA[21]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(21),
  I1 => cpi_lddata(21),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(21),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(21));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M_RNO_1[0]\: LUT6 
generic map(
  INIT => X"F0F0F0F08B0FAAAA"
)
port map (
  I0 => cpi_d_inst(10),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(63),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14_2\(77),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.TEMP_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8109\);
\GRLFPC20.WRDATA[26]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(26),
  I1 => cpi_lddata(26),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(26),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(26));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.NOTABORTWB_Z6648\: LUT6 
generic map(
  INIT => X"0F2F2F2F2F2F2F2F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(46),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14_2\(77),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\(5),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.OPREXCSHFT.UN3_OPREXC\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.NOTABORTWB\);
\GRLFPC20.R.I.EXC_RNIUP9M[5]\: LUT4 
generic map(
  INIT => X"007F"
)
port map (
  I0 => \GRLFPC20.R.I.EXC\(5),
  I1 => \GRLFPC20.R.I.V\,
  I2 => \GRLFPC20.COMB.V.I.EXEC_5\,
  I3 => \GRLFPC20.N_2000\,
  O => \GRLFPC20.N_3050\);
\GRLFPC20.WRDATA[60]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(28),
  I1 => cpi_lddata(28),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(60),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(28));
\GRLFPC20.WRDATA[57]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(25),
  I1 => cpi_lddata(25),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(57),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(25));
\GRLFPC20.WRDATA[28]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(28),
  I1 => cpi_lddata(28),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(28),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(28));
\GRLFPC20.WRDATA[31]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(31),
  I1 => cpi_lddata(31),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(31),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(31));
\GRLFPC20.WRDATA[30]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(30),
  I1 => cpi_lddata(30),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(30),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(30));
\GRLFPC20.WRDATA[0]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(0),
  I1 => cpi_lddata(0),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(0),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(0));
\GRLFPC20.WRDATA[1]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(1),
  I1 => cpi_lddata(1),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(1),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(1));
\GRLFPC20.WRDATA[2]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(2),
  I1 => cpi_lddata(2),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(2),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(2));
\GRLFPC20.WRDATA[3]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(3),
  I1 => cpi_lddata(3),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(3),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(3));
\GRLFPC20.WRDATA[4]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(4),
  I1 => cpi_lddata(4),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(4),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(4));
\GRLFPC20.WRDATA[5]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(5),
  I1 => cpi_lddata(5),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(5),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(5));
\GRLFPC20.WRDATA[6]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(6),
  I1 => cpi_lddata(6),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(6),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(6));
\GRLFPC20.WRDATA[7]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(7),
  I1 => cpi_lddata(7),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(7),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(7));
\GRLFPC20.WRDATA[8]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(8),
  I1 => cpi_lddata(8),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(8),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(8));
\GRLFPC20.WRDATA[9]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(9),
  I1 => cpi_lddata(9),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(9),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(9));
\GRLFPC20.WRDATA[10]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(10),
  I1 => cpi_lddata(10),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(10),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(10));
\GRLFPC20.WRDATA[11]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(11),
  I1 => cpi_lddata(11),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(11),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(11));
\GRLFPC20.WRDATA[12]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(12),
  I1 => cpi_lddata(12),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(12),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(12));
\GRLFPC20.WRDATA[13]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(13),
  I1 => cpi_lddata(13),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(13),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(13));
\GRLFPC20.WRDATA[14]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(14),
  I1 => cpi_lddata(14),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(14),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(14));
\GRLFPC20.WRDATA[15]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(15),
  I1 => cpi_lddata(15),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(15),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(15));
\GRLFPC20.WRDATA[16]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(16),
  I1 => cpi_lddata(16),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(16),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(16));
\GRLFPC20.WRDATA[17]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(17),
  I1 => cpi_lddata(17),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(17),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(17));
\GRLFPC20.WRDATA[18]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(18),
  I1 => cpi_lddata(18),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(18),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(18));
\GRLFPC20.WRDATA[19]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(19),
  I1 => cpi_lddata(19),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(19),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(19));
\GRLFPC20.WRDATA[20]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(20),
  I1 => cpi_lddata(20),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(20),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(20));
\GRLFPC20.WRDATA[22]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(22),
  I1 => cpi_lddata(22),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(22),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(22));
\GRLFPC20.WRDATA[23]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(23),
  I1 => cpi_lddata(23),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(23),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(23));
\GRLFPC20.WRDATA[24]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(24),
  I1 => cpi_lddata(24),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(24),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(24));
\GRLFPC20.WRDATA[25]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(25),
  I1 => cpi_lddata(25),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(25),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(25));
\GRLFPC20.WRDATA[27]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(27),
  I1 => cpi_lddata(27),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(27),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(27));
\GRLFPC20.WRDATA[29]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(29),
  I1 => cpi_lddata(29),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(29),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi2_wrdata(29));
\GRLFPC20.WRDATA[32]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(0),
  I1 => cpi_lddata(0),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(32),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(0));
\GRLFPC20.WRDATA[33]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(1),
  I1 => cpi_lddata(1),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(33),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(1));
\GRLFPC20.WRDATA[34]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(2),
  I1 => cpi_lddata(2),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(34),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(2));
\GRLFPC20.WRDATA[35]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(3),
  I1 => cpi_lddata(3),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(35),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(3));
\GRLFPC20.WRDATA[36]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(4),
  I1 => cpi_lddata(4),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(36),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(4));
\GRLFPC20.WRDATA[37]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(5),
  I1 => cpi_lddata(5),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(37),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(5));
\GRLFPC20.WRDATA[38]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(6),
  I1 => cpi_lddata(6),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(38),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(6));
\GRLFPC20.WRDATA[39]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(7),
  I1 => cpi_lddata(7),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(39),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(7));
\GRLFPC20.WRDATA[40]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(8),
  I1 => cpi_lddata(8),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(40),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(8));
\GRLFPC20.WRDATA[41]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(9),
  I1 => cpi_lddata(9),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(41),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(9));
\GRLFPC20.WRDATA[42]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(10),
  I1 => cpi_lddata(10),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(42),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(10));
\GRLFPC20.WRDATA[43]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(11),
  I1 => cpi_lddata(11),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(43),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(11));
\GRLFPC20.WRDATA[44]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(12),
  I1 => cpi_lddata(12),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(44),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(12));
\GRLFPC20.WRDATA[45]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(13),
  I1 => cpi_lddata(13),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(45),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(13));
\GRLFPC20.WRDATA[46]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(14),
  I1 => cpi_lddata(14),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(46),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(14));
\GRLFPC20.WRDATA[47]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(15),
  I1 => cpi_lddata(15),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(47),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(15));
\GRLFPC20.WRDATA[48]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(16),
  I1 => cpi_lddata(16),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(48),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(16));
\GRLFPC20.WRDATA[49]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(17),
  I1 => cpi_lddata(17),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(49),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(17));
\GRLFPC20.WRDATA[50]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(18),
  I1 => cpi_lddata(18),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(50),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(18));
\GRLFPC20.WRDATA[51]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(19),
  I1 => cpi_lddata(19),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(51),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(19));
\GRLFPC20.WRDATA[52]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(20),
  I1 => cpi_lddata(20),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(52),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(20));
\GRLFPC20.WRDATA[53]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(21),
  I1 => cpi_lddata(21),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(53),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(21));
\GRLFPC20.WRDATA[54]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(22),
  I1 => cpi_lddata(22),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(54),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(22));
\GRLFPC20.WRDATA[55]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(23),
  I1 => cpi_lddata(23),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(55),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(23));
\GRLFPC20.WRDATA[56]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(24),
  I1 => cpi_lddata(24),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(56),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(24));
\GRLFPC20.WRDATA[58]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(26),
  I1 => cpi_lddata(26),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(58),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(26));
\GRLFPC20.WRDATA[59]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(27),
  I1 => cpi_lddata(27),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(59),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(27));
\GRLFPC20.WRDATA[61]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(29),
  I1 => cpi_lddata(29),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(61),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(29));
\GRLFPC20.WRDATA[62]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(30),
  I1 => cpi_lddata(30),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.WRDATA_4\(62),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(30));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_154_I_X2\: LUT5_L 
generic map(
  INIT => X"87878877"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\(35),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(35),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_841_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_106_I_X2\: LUT5_L 
generic map(
  INIT => X"87878877"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\(38),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(38),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_838_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_74_I_X2\: LUT5_L 
generic map(
  INIT => X"87878877"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(56),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_836_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M_RNO_0[0]\: LUT5 
generic map(
  INIT => X"CC0ACCFA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(60),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_10\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[7]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1272\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10157_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1748\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(7),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2\(7),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[49]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1650\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2125\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_1\(49),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_2\(49),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_2\(49),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(49));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[4]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFF8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2602\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1580\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_0\(4),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(4),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1710\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_3\(4),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[55]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7\(55),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_1\(55),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(55),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2\(55),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8\(55),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9\(55),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(55));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[27]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2831\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12248\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(27),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7\(27),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(27),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_0\(27),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(27));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[25]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF08"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_7_1\(25),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9968_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1536_I\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9720\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_0\(25),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(25),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(25));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[18]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9605\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9601\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(18),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3\(18),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5\(18),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(18),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(18));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I[31]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9385\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_6_0\(31),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_2\(31),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_6_1\(31),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_7_0\(31),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_0_1\(31),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(31));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[57]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10605\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10678\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_1\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4\(57),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(57),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_13\(57),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[19]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_0\(19),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_1\(19),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8\(19),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7\(19),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(19),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[6]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_1\(6),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_0\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2140\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4\(6),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(6),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7\(6),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[0]\: LUT5_L 
generic map(
  INIT => X"FFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9445\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1039\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9453\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(0),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[59]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1229\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1169\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7\(59),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5\(59),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(59),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(59));
\GRLFPC20.RS1_1_0[1]\: LUT6 
generic map(
  INIT => X"FFFF2020FFFF3300"
)
port map (
  I0 => cpi_d_inst(15),
  I1 => cpi_dbg_enable,
  I2 => \GRLFPC20.N_1583\,
  I3 => \GRLFPC20.R.A.RS1\(1),
  I4 => \GRLFPC20.RS1_1_0_0\(1),
  I5 => holdn,
  O => RFI2_RD1ADDR_16);
\GRLFPC20.RS1_1_0[2]\: LUT6 
generic map(
  INIT => X"FFFF2020FFFF3300"
)
port map (
  I0 => cpi_d_inst(16),
  I1 => cpi_dbg_enable,
  I2 => \GRLFPC20.N_1583\,
  I3 => \GRLFPC20.R.A.RS1\(2),
  I4 => \GRLFPC20.RS1_1_0_0\(2),
  I5 => holdn,
  O => RFI2_RD1ADDR_17);
\GRLFPC20.RS1_1_0[3]\: LUT6 
generic map(
  INIT => X"FFFF2020FFFF3300"
)
port map (
  I0 => cpi_d_inst(17),
  I1 => cpi_dbg_enable,
  I2 => \GRLFPC20.N_1583\,
  I3 => \GRLFPC20.R.A.RS1\(3),
  I4 => \GRLFPC20.RS1_1_0_0\(3),
  I5 => holdn,
  O => RFI2_RD1ADDR_18);
\GRLFPC20.RS1_1_0[4]\: LUT6 
generic map(
  INIT => X"FFFF2020FFFF3300"
)
port map (
  I0 => cpi_d_inst(18),
  I1 => cpi_dbg_enable,
  I2 => \GRLFPC20.N_1583\,
  I3 => \GRLFPC20.R.A.RS1\(4),
  I4 => \GRLFPC20.RS1_1_0_0\(4),
  I5 => holdn,
  O => RFI2_RD1ADDR_19);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[12]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFA8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10157_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2774\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1283\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2337\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1661\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3\(12),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(12));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[5]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_982\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_0\(5),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_966\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3\(5),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_4\(5),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_1\(5),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[50]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFF8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10157_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1342\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3\(50),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2151\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2\(50),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1\(50),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(50));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_11[52]_Z6735\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFF8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2605\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10246_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(52),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7_1\(52),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4\(52),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5\(52),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_11\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2_2[60]_Z6736\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFF8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10157_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1282\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_7\(60),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2_0\(60),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2_1\(60),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_5\(60),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2_2\(60));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_17[75]\: LUT6_L 
generic map(
  INIT => X"0F87F087F087F087"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(9),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(48),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(52),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\(5),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\(3),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8821\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"F20D20DF0DF2DF20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(318),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(55),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.CIN_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.SI_6\(51),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.SI_64\(49));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"F20D20DF0DF2DF20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(333),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(40),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.CIN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.SI_21\(36),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.SI_79\(34));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"2DD2D22DD22D2DD2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(331),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(42),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.CIN_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.CIN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.SI_78\(35));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"F20D20DF0DF2DF20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(328),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(45),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.CIN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.CIN_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.SI_16\(41),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.SI_74\(39));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"F20D20DF0DF2DF20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(326),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(47),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.CIN_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.SI_14\(43),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.SI_72\(41));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"2DD2D22DD22D2DD2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(324),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.CIN_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.CIN_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.SI_71\(42));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"F20D20DF0DF2DF20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(324),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.CIN_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.CIN_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.SI_12\(45),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.SI_70\(43));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"AC0053FF53FFAC00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.UN195_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.UN198_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10.Z_C1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.SI_10\(47),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.SI_68\(45));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"2DD2D22DD22D2DD2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(318),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(55),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.CIN_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.SI_65\(48));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"2DD2D22DD22D2DD2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(346),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(27),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.CIN_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.SI_93\(20));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"AC0053FF53FFAC00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.UN252_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.UN255_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_C1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.SI_29\(28),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.SI_87\(26));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"2DD2D22DD22D2DD2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(338),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(35),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.CIN_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.CIN_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.SI_85\(28));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"F20D20DF0DF2DF20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(338),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(35),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.CIN_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.CIN_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.SI_26\(31),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.SI_84\(29));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"2DD2D22DD22D2DD2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(333),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(40),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.CIN_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.SI_80\(33));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"0DF2DF20F20D20DF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(357),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(16),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_541\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.CIN_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.SI_45\(12),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.SI_103\(10));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"0DF2DF20F20D20DF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(355),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(18),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_548\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.SI_43\(14),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.SI_101\(12));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"D22D2DD22DD2D22D"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(353),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(20),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_550\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.CIN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.SI_100\(13));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"F20D20DF0DF2DF20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(351),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(22),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_559\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.CIN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.SI_39\(18),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.SI_97\(16));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39.Z_AC0_1_Z6756\: LUT6 
generic map(
  INIT => X"00F20020F2002000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(351),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(22),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_559\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.CIN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.SI_39\(18),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39.Z_AC0_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"F20D20DF0DF2DF20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(349),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(24),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.CIN_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.CIN_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.SI_37\(20),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.SI_95\(18));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51.Z_AC0_1_Z6758\: LUT6 
generic map(
  INIT => X"F200200000F20020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(363),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(10),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_515\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.SI_51\(6),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51.Z_AC0_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"AC0053FF53FFAC00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_811_I\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_812_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50.Z_C1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.SI_50\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.SI_108\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"0DF2DF20F20D20DF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(359),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(14),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_523\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.CIN_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.SI_47\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.SI_105\(8));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI3CFC3_0[368]\: LUT6 
generic map(
  INIT => X"F20D20DF0DF2DF20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(368),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(5),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.SI_56\(1),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SBLSBS_1\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL_AXBXC1\: LUT3 
generic map(
  INIT => X"A6"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  O => N_4325);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[38]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFF4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_775\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2772\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2235\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_969\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_972\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1776\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(38));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[53]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10310\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10292\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10309\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4\(53),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(53),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9\(53),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(53));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[34]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFF8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_1_0\(36),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9957\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9964\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2\(34),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(34),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(34),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRLOI\(34));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_RNID0RF2\: LUT6_L 
generic map(
  INIT => X"2DD2D22DD22D2DD2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(368),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(5),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO0_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SBLSBS_2\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIQNCS3[368]\: LUT6 
generic map(
  INIT => X"2DD2D22DD22D2DD2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(368),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(5),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.CIN_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN16_NOTPROP_2336_0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO0_0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN16_NOTPROP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_58_0_A2[56]\: LUT6 
generic map(
  INIT => X"39FFC600C60039FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2963_I\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12044\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0_0[0]\: LUT6 
generic map(
  INIT => X"EAEAEAEAEEAAEEEE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0_0_0\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0_0_A2_0\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M13\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M12\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_I_I_A2_0_O2_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_SM12\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0_0_O2[2]\: LUT6 
generic map(
  INIT => X"EAEAEAEAEEAAEEEE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0_0_O2_0\(2),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0_0_A2_0\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M13\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M12\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_I_I_A2_0_O2_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_SM12\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_I_A2_RNIUKD71[0]\: LUT5_L 
generic map(
  INIT => X"000000A2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(38),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(39),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(40),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1186\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1101\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_593_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[45]_Z6772\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(186),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(45));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[51]_Z6773\: LUT6 
generic map(
  INIT => X"000000CC00F0AA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(180),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(51));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[52]_Z6774\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(179),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[44]_Z6775\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(187),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(44));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN3_NOTRESETORUNIMP_Z6776\: LUT4 
generic map(
  INIT => X"050D"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(66),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(67),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.ENTRYPOINT\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN3_NOTRESETORUNIMP\);
\GRLFPC20.COMB.SEQERR.UN7_OP\: LUT4 
generic map(
  INIT => X"FF80"
)
port map (
  I0 => cpi_d_inst(30),
  I1 => cpi_d_inst(31),
  I2 => \GRLFPC20.N_1142\,
  I3 => \GRLFPC20.N_1583\,
  O => \GRLFPC20.N_1138\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[5]_Z6778\: LUT6 
generic map(
  INIT => X"000000CC00F0AA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(226),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[22]_Z6779\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(209),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(22));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[12]_Z6780\: LUT6 
generic map(
  INIT => X"000000CC00F0AA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(219),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(12));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[22]_Z6781\: LUT6 
generic map(
  INIT => X"F7B3D591E6A2C480"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8233\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8234\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8235\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8236\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(22));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[23]_Z6782\: LUT6 
generic map(
  INIT => X"F7B3D591E6A2C480"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8232\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8233\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8234\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8235\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(23));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[24]_Z6783\: LUT6 
generic map(
  INIT => X"F7B3D591E6A2C480"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8231\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8232\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8233\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8234\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(24));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[25]_Z6784\: LUT6 
generic map(
  INIT => X"F7B3D591E6A2C480"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8230\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8231\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8232\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8233\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(25));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[21]_Z6785\: LUT6 
generic map(
  INIT => X"FE76BA32DC549810"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8237\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8234\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8235\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8236\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(21));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[56]_Z6786\: LUT6 
generic map(
  INIT => X"F7B3E6A2D591C480"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8199\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8200\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8202\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8201\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(56));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[57]_Z6787\: LUT6 
generic map(
  INIT => X"F7B3D591E6A2C480"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8198\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8199\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8200\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8201\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[12]_Z6788\: LUT6 
generic map(
  INIT => X"FE76BA32DC549810"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8246\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8243\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8244\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8245\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(12));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[55]_Z6789\: LUT6 
generic map(
  INIT => X"F7D5E6C4B391A280"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8200\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8202\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8203\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8201\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(55));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[54]_Z6790\: LUT6 
generic map(
  INIT => X"FEBADC9876325410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8204\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8202\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8203\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8201\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[1]_Z6791\: LUT5 
generic map(
  INIT => X"FF7F8000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(56),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(57),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[2]_Z6792\: LUT6 
generic map(
  INIT => X"FF7FBF3FC0408000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(55),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(56),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(57),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[43]_Z6793\: LUT6 
generic map(
  INIT => X"000000CC00F0AA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(188),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(43));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[27]_Z6794\: LUT6 
generic map(
  INIT => X"000000CC00F0AA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(204),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(27));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[2]_Z6795\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(229),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[13]_Z6796\: LUT6 
generic map(
  INIT => X"F7B3D591E6A2C480"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8242\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8243\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8244\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8245\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(13));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[14]_Z6797\: LUT6 
generic map(
  INIT => X"F7B3D591E6A2C480"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8241\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8242\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8243\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8244\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(14));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[45]_Z6798\: LUT6 
generic map(
  INIT => X"F7B3D591E6A2C480"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8210\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8211\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8212\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8213\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(45));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[44]_Z6799\: LUT6 
generic map(
  INIT => X"F7E6B3A2D5C49180"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8211\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8214\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8212\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8213\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(44));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[43]_Z6800\: LUT6 
generic map(
  INIT => X"FDEC7564B9A83120"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8214\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8215\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8212\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8213\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(43));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[20]_Z6801\: LUT6 
generic map(
  INIT => X"FDEC7564B9A83120"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8237\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8238\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8235\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8236\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(20));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[3]_Z6802\: LUT6 
generic map(
  INIT => X"55154000FFBFEAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(55),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(57),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[55]_Z6803\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(176),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(55));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[54]_Z6804\: LUT6 
generic map(
  INIT => X"000000CC00F0AA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(177),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[53]_Z6805\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(178),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(53));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[50]_Z6806\: LUT6 
generic map(
  INIT => X"000000CC00F0AA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(181),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(50));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[49]_Z6807\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(182),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(49));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[48]_Z6808\: LUT6 
generic map(
  INIT => X"000000CC00F0AA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(183),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(48));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[47]_Z6809\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(184),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[46]_Z6810\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(185),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(46));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[42]_Z6811\: LUT6 
generic map(
  INIT => X"000000CC00F0AA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(189),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(42));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[41]_Z6812\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(190),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(41));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[40]_Z6813\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(191),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(40));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[39]_Z6814\: LUT6 
generic map(
  INIT => X"000000CC00F0AA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(192),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(39));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[32]_Z6815\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(199),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(32));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[31]_Z6816\: LUT6 
generic map(
  INIT => X"000000CC00F0AA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(200),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(31));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[29]_Z6817\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(202),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(29));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[28]_Z6818\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(203),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(28));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[21]_Z6819\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(210),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(21));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[20]_Z6820\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(211),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(20));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[19]_Z6821\: LUT6 
generic map(
  INIT => X"000000CC00F0AA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(212),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[18]_Z6822\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(213),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(18));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[17]_Z6823\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(214),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(17));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[16]_Z6824\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(215),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(16));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[15]_Z6825\: LUT6 
generic map(
  INIT => X"000000CC00F0AA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(216),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(15));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[14]_Z6826\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(217),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(14));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[13]_Z6827\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(218),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(13));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[11]_Z6828\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(220),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[10]_Z6829\: LUT6 
generic map(
  INIT => X"000000CC00F0AA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(221),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(10));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[9]_Z6830\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(222),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(9));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[8]_Z6831\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(223),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(8));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[7]_Z6832\: LUT6 
generic map(
  INIT => X"000000CC00F0AA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(224),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[6]_Z6833\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(225),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[4]_Z6834\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(227),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[3]_Z6835\: LUT6 
generic map(
  INIT => X"000000CC00F0AA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(228),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[42]\: LUT5_L 
generic map(
  INIT => X"FFFFFFF8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2608\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10157_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2219\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1\(42),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1653\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(42));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[44]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF10"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_254\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10157_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(44),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0\(44),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1748\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(44));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[30]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFEAC0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12195\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1335\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1234\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2818\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_866\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_1\(30),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRLOI\(30));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[3]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0504"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_715\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2605\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2608\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2559\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2\(3),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[26]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF10"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_289\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2600\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1593\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0\(26),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1\(26),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(26));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[28]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2695\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_291_I\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_0\(28),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_1\(28),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2\(28),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(28));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[13]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF10"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9610_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9785_1_I_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1169\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3\(13),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5\(13),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4\(13),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(13));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[36]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10016\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9549_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9667_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(36),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3\(36),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8\(36),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(36));
\GRLFPC20.RS1V_0_SQMUXA_1_Z6844\: LUT6 
generic map(
  INIT => X"1010100000000000"
)
port map (
  I0 => cpi_d_inst(19),
  I1 => cpi_d_inst(20),
  I2 => cpi_d_inst(23),
  I3 => \GRLFPC20.N_3081\,
  I4 => \GRLFPC20.N_3082\,
  I5 => \GRLFPC20.N_3109\,
  O => \GRLFPC20.RS1V_0_SQMUXA_1\);
\GRLFPC20.COMB.RS2D_1_IV\: LUT6 
generic map(
  INIT => X"FEFAFAFAFCF0F0F0"
)
port map (
  I0 => \GRLFPC20.N_925\,
  I1 => \GRLFPC20.N_3083_1\,
  I2 => \GRLFPC20.N_3106\,
  I3 => \GRLFPC20.N_3120\,
  I4 => \GRLFPC20.N_3129\,
  I5 => \GRLFPC20.COMB.FPDECODE.RS1D5\,
  O => \GRLFPC20.COMB.RS2D_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15[16]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFF1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_135\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_765\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2233\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2156\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15_0_0\(16),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15_1\(16),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(16));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14[77]_Z6847\: LUT6 
generic map(
  INIT => X"0020202020202020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(46),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14_2\(77),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\(5),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.OPREXCSHFT.UN3_OPREXC\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14\(77));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6[25]_Z6848\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF02"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1132_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10790\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_406\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9716\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(25),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2\(25),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(25));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6[32]_Z6849\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFFF80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9863_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_991_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1041\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0\(32),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(32));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_7[11]_Z6850\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFFF20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_717\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10626_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9323\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_0\(11),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_7_0\(11),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_7\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_13[57]_Z6851\: LUT5_L 
generic map(
  INIT => X"FFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10609\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9\(57),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(57),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_11\(57),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_13\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6[33]_Z6852\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFFF10"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9887_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2594\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2734\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(33),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_1\(33),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(33));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1[51]_Z6853\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2590\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_921\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9394_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10157\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1654\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_0\(51),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(51));
\GRLFPC20.COMB.V.FSR.CEXC_1_IV_0[2]_Z6854\: LUT5 
generic map(
  INIT => X"B8888888"
)
port map (
  I0 => cpi_dbg_data(2),
  I1 => \GRLFPC20.N_1704\,
  I2 => \GRLFPC20.R.I.EXC\(2),
  I3 => \GRLFPC20.R.FSR.TEM\(2),
  I4 => \GRLFPC20.N_2000\,
  O => \GRLFPC20.COMB.V.FSR.CEXC_1_IV_0\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_18[74]_Z6855\: LUT6_L 
generic map(
  INIT => X"008AAAAAAAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(62),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CONDMUXMULXFF.UN5_NOTSQRTLFTCC\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_WQSTSETS\(0),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_18\(74));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_3_RNI5S3U_0\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(312),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(370),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7498_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIP5M92[24]\: LUT6 
generic map(
  INIT => X"ACFF00FF5300FF00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SALSBS_2\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN10_NOTPROP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIP5M92_0[24]\: LUT6 
generic map(
  INIT => X"5300FF0000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SALSBS_2\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN12_GEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1_Z6859\: LUT4 
generic map(
  INIT => X"00FB"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(71),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(75),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIAML61_0[311]\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(311),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(369),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO0_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6.Z_C1_Z6861\: LUT4 
generic map(
  INIT => X"F220"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(318),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(55),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5.Z_C1_Z6862\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(259),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(317),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_C1_Z6863\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(274),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(332),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.CIN_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19.Z_C1_Z6864\: LUT4 
generic map(
  INIT => X"F220"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(331),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(42),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.CIN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18.Z_C1_Z6865\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(272),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(330),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.CIN_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_C1_Z6866\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(271),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(329),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_AXB1_Z6867\: LUT5 
generic map(
  INIT => X"D22D2DD2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(328),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(45),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.CIN_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.CIN_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_AXB1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_C1_Z6868\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(269),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(327),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.CIN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_C1_Z6869\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(267),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(325),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.CIN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11.Z_C1_Z6870\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(265),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(323),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10.Z_C1_Z6871\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(264),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(322),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.CIN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9.Z_C1_Z6872\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(263),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(321),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8.Z_C1_Z6873\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(262),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(320),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7.Z_C1_Z6874\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(261),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(319),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36.Z_C1_Z6875\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(290),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(348),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35.Z_C1_Z6876\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(289),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(347),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_C1_Z6877\: LUT4 
generic map(
  INIT => X"F220"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(346),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(27),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33.Z_C1_Z6878\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(287),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(345),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.CIN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_C1_Z6879\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(286),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(344),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31.Z_C1_Z6880\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(285),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(343),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_C1_Z6881\: LUT4 
generic map(
  INIT => X"F220"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(342),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(31),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.CIN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_C1_Z6882\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(283),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(341),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.CIN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28.Z_C1_Z6883\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(282),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(340),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.CIN_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27.Z_C1_Z6884\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(281),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(339),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.CIN_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26.Z_AXB1_Z6885\: LUT6 
generic map(
  INIT => X"3A0AC5F5C5F53A0A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(279),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_AXB0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26.Z_AXB1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_C1_Z6886\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(279),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(337),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24.Z_C1_Z6887\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(278),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(336),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_C1_Z6888\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(277),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(335),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.CIN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_AXB1_Z6889\: LUT6 
generic map(
  INIT => X"C3A5FFFF3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.SI_23\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_AXB1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_AC0_2_Z6890\: LUT6 
generic map(
  INIT => X"3C5A000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.SI_23\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_AC0_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22.Z_C1_Z6891\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(276),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(334),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44.Z_C1_Z6892\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(298),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(356),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_C1_Z6893\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(296),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(354),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38.Z_C1_Z6894\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(292),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(350),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50.Z_C1_Z6895\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(304),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(362),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.CIN_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49.Z_C1_Z6896\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(303),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(361),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_C1_Z6897\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(300),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(358),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_AXB1_Z6898\: LUT5 
generic map(
  INIT => X"2DD2D22D"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(357),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(16),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_537\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_AXB1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55.Z_C1_Z6899\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(309),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(367),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53.Z_C1_Z6900\: LUT6 
generic map(
  INIT => X"0FEE00EE00880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(307),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(365),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[37]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2590\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1169\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(37),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0\(37),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_782\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(37));
\GRLFPC20.RS1D_CNST.M10\: LUT5 
generic map(
  INIT => X"20000000"
)
port map (
  I0 => cpi_d_inst(21),
  I1 => cpi_d_inst(22),
  I2 => cpi_d_inst(24),
  I3 => cpi_d_inst(31),
  I4 => \GRLFPC20.RS1D_CNST.N_7\,
  O => \GRLFPC20.RS1D_CNST\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[61]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF8C"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10895\,
  I1 => N_3105_TZ,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_222\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10891\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(61),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5\(61),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(61));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_I_26\: LUT6 
generic map(
  INIT => X"8124184200000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(6),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(7),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12036\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_N_11\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_0_Z6905\: LUT6_L 
generic map(
  INIT => X"FF22F020F020F020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_2_I\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_6\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR_0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR_1\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[23]_Z6906\: LUT6 
generic map(
  INIT => X"000000CC00F0AA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(208),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(23));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[24]_Z6907\: LUT6 
generic map(
  INIT => X"000000CC00F0AA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(207),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(24));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[30]_Z6908\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(201),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(30));
\GRLFPC20.COMB.V.I.RES_1[63]_Z6909\: LUT6_L 
generic map(
  INIT => X"5F500F005C5C0C0C"
)
port map (
  I0 => cpi_a_inst(8),
  I1 => \GRLFPC20.R.I.RES\(63),
  I2 => \GRLFPC20.N_1858\,
  I3 => \GRLFPC20.FPO.SIGN\,
  I4 => \GRLFPC20.COMB.UN15_HOLDN\,
  I5 => \GRLFPC20.N_2102\,
  LO => \GRLFPC20.COMB.V.I.RES_1\(63));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_39_1[0]\: LUT6 
generic map(
  INIT => X"3C3CFF005A5AFF00"
)
port map (
  I0 => rfo1_data2(31),
  I1 => rfo2_data2(31),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(0),
  I3 => \GRLFPC20.FPO.SIGN\,
  I4 => \GRLFPC20.FPI.LDOP\,
  I5 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9257\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[25]_Z6911\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(206),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(25));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1[26]_Z6912\: LUT6 
generic map(
  INIT => X"000000F000CCAA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(205),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(26));
\GRLFPC20.COMB.UN1_MEXC_1_0_LUT6_2_RNIC2242\: LUT6 
generic map(
  INIT => X"0002000000000000"
)
port map (
  I0 => \GRLFPC20.R.I.V\,
  I1 => \GRLFPC20.N_1306\,
  I2 => \GRLFPC20.N_1307\,
  I3 => \GRLFPC20.N_1310\,
  I4 => \GRLFPC20.COMB.UN1_MEXC_1_0\,
  I5 => \GRLFPC20.COMB.V.I.EXEC_5\,
  O => \GRLFPC20.N_2146\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_0_YY[2]\: LUT5 
generic map(
  INIT => X"0F0F2D87"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => N_6675);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_0_YY[3]\: LUT5 
generic map(
  INIT => X"0F0F2D87"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => N_6683);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_0_YY[4]\: LUT5 
generic map(
  INIT => X"0F0F2D87"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => N_6691);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[41]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFF808080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9394_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9861_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2608\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10157_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1282\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1\(41),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(41));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[1]\: LUT3_L 
generic map(
  INIT => X"FE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2831\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2559\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1726\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_O2[24]\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFFF20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1536_I\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_830\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2608\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1187\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1039\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_O2_0\(24),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1775\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_0_A2[2]\: LUT5_L 
generic map(
  INIT => X"00000020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(38),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(39),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(40),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1186\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1101\,
  LO => \GRLFPC20.FPO.EXC\(2));
\GRLFPC20.UN1_FPOP7_0_A3\: LUT5 
generic map(
  INIT => X"10000000"
)
port map (
  I0 => cpi_d_inst(8),
  I1 => cpi_d_inst(13),
  I2 => \GRLFPC20.N_3079\,
  I3 => \GRLFPC20.N_3128\,
  I4 => \GRLFPC20.N_3129\,
  O => \GRLFPC20.N_3106\);
\GRLFPC20.MOV_5_SQMUXA_0_A3\: LUT6_L 
generic map(
  INIT => X"0007000000000000"
)
port map (
  I0 => cpi_d_inst(7),
  I1 => cpi_d_inst(8),
  I2 => cpi_d_inst(10),
  I3 => cpi_d_inst(11),
  I4 => \GRLFPC20.N_3127\,
  I5 => \GRLFPC20.N_3129\,
  LO => \GRLFPC20.N_865\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0[35]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFECA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2697\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10223_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2591\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10626_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2255\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(35),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(35));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[23]\: LUT5_L 
generic map(
  INIT => X"FFFFEAC0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9453_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2594\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2608\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10157_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2\(23),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(23));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_1[30]_Z6925\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFF0C8C0C"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2337_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_85\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9861_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_789\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0\(30),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_1\(30));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8[36]_Z6926\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF08"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_15_1\(36),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_830\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10035\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2730\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0\(36),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8\(36));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6[27]_Z6927\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFFF10"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10006\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12021_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9\(27),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0\(27),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_0\(27),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(27));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_3[4]_Z6928\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFEAC0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_830\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1562\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_157_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2774\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10699\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2\(4),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_3\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_4[5]_Z6929\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFFF10"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_234\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1336\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(5),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1\(5),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1592\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_4\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2[50]_Z6930\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFF888"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_134_I\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_777\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_995_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10943\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2206\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0\(50),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2\(50));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2[7]_Z6931\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFECCCA000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10592_I\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9601_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10025_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2600\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2505_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_0\(7),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5[59]_Z6932\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFF888"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10724\,
  I1 => N_3154_TZ,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_314_I\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2701\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10751\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(59),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5\(59));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6[59]_Z6933\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF04"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_52\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10765_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_906\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10748\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0\(59),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_0\(59),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(59));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8[32]_Z6934\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF08"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9390_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9911_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_304\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9846\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2125\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0\(32),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8\(32));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3[12]_Z6935\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2475\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_965\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9860\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_967\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_966\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1\(12),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3\(12));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_7[47]_Z6936\: LUT6 
generic map(
  INIT => X"FFFFFFFFC0C0EAC0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2693\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_6_0\(47),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10943\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_765\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_0\(47),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_7\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2_1[47]_Z6937\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10834\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10082\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_1_0\(47),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_6_1\(47),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_4\(47),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_6_0\(47),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2_1\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2_1[11]_Z6938\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFFF80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9667_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9492_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9738_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_4_0\(11),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_3\(11),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_1_1\(11),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2_1\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6[6]_Z6939\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFFFF8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_7_0\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2724\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9974\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9497\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(6),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(6),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_1[17]_Z6940\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFFFF4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2831\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_981\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2159\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1592\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_0\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_1\(17));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9[33]_Z6941\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9925_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_59\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9600_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9922\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_0\(33),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8\(33),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9\(33));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7[58]_Z6942\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF0C0E"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10696_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10661\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_409\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9451\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7_1\(58),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7\(58));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8[58]_Z6943\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A30_23_0\(58),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9969_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_314_I\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10699\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0\(58),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8_2\(58),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8\(58));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7[54]_Z6944\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFFF08"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1232\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12131\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10365\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_0\(54),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7_1\(54),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_6_2[60]_Z6945\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFFF20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10293_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_428\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9652_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_1_0\(60),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_0\(60),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_4\(60),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_6_2\(60));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_2[49]_Z6946\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9492_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10157_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2151\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_0\(49),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_1\(49),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_2\(49));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_7_0[56]_Z6947\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFF2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_7_TZ\(56),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1006\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10524\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_3\(56),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_1\(56),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_7_0\(56));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_8[56]_Z6948\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFF400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_759\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9408_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9453_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_6\(56),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2\(56),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_8\(56));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_1[51]_Z6949\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF1110"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_766\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2605\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2608\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_5_0\(51),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_5_1\(51),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_1\(51));
\GRLFPC20.V.I.V_3_SQMUXA_0_Z6950\: LUT5 
generic map(
  INIT => X"0000000B"
)
port map (
  I0 => \GRLFPC20.N_1295\,
  I1 => \GRLFPC20.R.X.SEQERR\,
  I2 => \GRLFPC20.N_1858\,
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.N_2000\,
  O => \GRLFPC20.V.I.V_3_SQMUXA_0\);
\GRLFPC20.R.I.EXEC_RNO_0\: LUT5 
generic map(
  INIT => X"FFFFD5FF"
)
port map (
  I0 => rst,
  I1 => \GRLFPC20.R.A.MOV\,
  I2 => \GRLFPC20.N_2931_1\,
  I3 => \GRLFPC20.COMB.V.I.EXEC_5\,
  I4 => \GRLFPC20.N_2000\,
  O => \GRLFPC20.COMB.V.I.EXEC_18_0_29_I_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[32]_Z6952\: LUT5 
generic map(
  INIT => X"0053FF53"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(27),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(31),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8223\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(32));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[34]_Z6953\: LUT5 
generic map(
  INIT => X"530053FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(23),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(27),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8223\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(34));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_3_RNI5S3U\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(312),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(370),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SALSBS_2\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[23]\: LUT5 
generic map(
  INIT => X"FACC0ACC"
)
port map (
  I0 => rfo2_data2(31),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(139),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  I4 => \GRLFPC20.FPI.OP2\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7894\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[7]_Z6956\: LUT6 
generic map(
  INIT => X"084C2A6E195D3B7F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(50),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(54),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(52),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(56),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[9]_Z6957\: LUT6 
generic map(
  INIT => X"02138A9B4657CEDF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(50),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(54),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(48),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(52),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(9));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[11]_Z6958\: LUT6 
generic map(
  INIT => X"40704C7C43734F7F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(46),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(50),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(48),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(52),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[17]_Z6959\: LUT5 
generic map(
  INIT => X"0053FF53"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(42),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(46),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8238\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(17));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[18]_Z6960\: LUT5 
generic map(
  INIT => X"0053FF53"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(41),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8237\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(18));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[26]_Z6961\: LUT5 
generic map(
  INIT => X"350035FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(35),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(31),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8231\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(26));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[28]_Z6962\: LUT5 
generic map(
  INIT => X"0035FF35"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(35),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(31),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8227\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(28));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[30]_Z6963\: LUT5 
generic map(
  INIT => X"530053FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(27),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(31),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8227\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(30));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[38]_Z6964\: LUT5 
generic map(
  INIT => X"530053FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(19),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(23),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8219\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(38));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[40]_Z6965\: LUT5 
generic map(
  INIT => X"0053FF53"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(19),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(23),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8215\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(40));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[10]_Z6966\: LUT6 
generic map(
  INIT => X"024613578ACE9BDF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(51),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(53),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(47),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(10));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[8]_Z6967\: LUT6 
generic map(
  INIT => X"082A4C6E193B5D7F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(51),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(53),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(55),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(8));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[6]_Z6968\: LUT6 
generic map(
  INIT => X"082A4C6E193B5D7F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(51),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(53),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(55),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(57),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[4]_Z6969\: LUT5 
generic map(
  INIT => X"082A5D7F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(53),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(55),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(57),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[16]_Z6970\: LUT6 
generic map(
  INIT => X"550F3300550F33FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(41),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(43),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(45),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(47),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(16));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[14]_Z6971\: LUT6 
generic map(
  INIT => X"5030503F5F305F3F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(43),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(49),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(47),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(14));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[12]\: LUT5 
generic map(
  INIT => X"FACA3A0A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(128),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.FPI.OP2\(42),
  I4 => \GRLFPC20.FPI.OP2\(45),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7905\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0[35]_Z6973\: LUT5 
generic map(
  INIT => X"CCCCCAAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(196),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(35));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0[34]_Z6974\: LUT5 
generic map(
  INIT => X"CCCCCAAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(197),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(34));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[15]_Z6975\: LUT6 
generic map(
  INIT => X"550F3300550F33FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(42),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(44),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(46),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(48),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(15));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[3]_Z6976\: LUT5 
generic map(
  INIT => X"082A5D7F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(54),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(56),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(57),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[5]_Z6977\: LUT6 
generic map(
  INIT => X"028A46CE139B57DF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(54),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(52),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(56),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(57),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(5));
\GRLFPC20.COMB.V.E.STDATA_1[22]_Z6978\: LUT5_L 
generic map(
  INIT => X"CACFCAC0"
)
port map (
  I0 => \GRLFPC20.R.FSR.NONSTD\,
  I1 => \GRLFPC20.N_2361\,
  I2 => \GRLFPC20.R.A.AFQ\,
  I3 => \GRLFPC20.R.A.AFSR\,
  I4 => \GRLFPC20.FPI.OP1\(54),
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(22));
\GRLFPC20.COMB.V.E.STDATA_1[0]_Z6979\: LUT6_L 
generic map(
  INIT => X"44F044FF44F04400"
)
port map (
  I0 => \GRLFPC20.COMB.V.E.STDATA2\,
  I1 => \GRLFPC20.R.I.INST\(0),
  I2 => \GRLFPC20.R.FSR.CEXC\(0),
  I3 => \GRLFPC20.R.A.AFQ\,
  I4 => \GRLFPC20.R.A.AFSR\,
  I5 => \GRLFPC20.FPI.OP1\(32),
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(0));
\GRLFPC20.COMB.V.E.STDATA_1[1]_Z6980\: LUT6_L 
generic map(
  INIT => X"44F044FF44F04400"
)
port map (
  I0 => \GRLFPC20.COMB.V.E.STDATA2\,
  I1 => \GRLFPC20.R.I.INST\(1),
  I2 => \GRLFPC20.R.FSR.CEXC\(1),
  I3 => \GRLFPC20.R.A.AFQ\,
  I4 => \GRLFPC20.R.A.AFSR\,
  I5 => \GRLFPC20.FPI.OP1\(33),
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(1));
\GRLFPC20.COMB.V.E.STDATA_1[6]_Z6981\: LUT5_L 
generic map(
  INIT => X"CACFCAC0"
)
port map (
  I0 => \GRLFPC20.R.FSR.AEXC\(1),
  I1 => \GRLFPC20.N_2345\,
  I2 => \GRLFPC20.R.A.AFQ\,
  I3 => \GRLFPC20.R.A.AFSR\,
  I4 => \GRLFPC20.FPI.OP1\(38),
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(6));
\GRLFPC20.COMB.V.E.STDATA_1[8]_Z6982\: LUT5_L 
generic map(
  INIT => X"CACFCAC0"
)
port map (
  I0 => \GRLFPC20.R.FSR.AEXC\(3),
  I1 => \GRLFPC20.N_2347\,
  I2 => \GRLFPC20.R.A.AFQ\,
  I3 => \GRLFPC20.R.A.AFSR\,
  I4 => \GRLFPC20.FPI.OP1\(40),
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(8));
\GRLFPC20.COMB.V.E.STDATA_1[15]_Z6983\: LUT5_L 
generic map(
  INIT => X"CACFCAC0"
)
port map (
  I0 => \GRLFPC20.R.FSR.FTT\(1),
  I1 => \GRLFPC20.N_2354\,
  I2 => \GRLFPC20.R.A.AFQ\,
  I3 => \GRLFPC20.R.A.AFSR\,
  I4 => \GRLFPC20.FPI.OP1\(47),
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(15));
\GRLFPC20.COMB.V.FSR.TEM_1[4]_Z6984\: LUT6_L 
generic map(
  INIT => X"A0C0A0C0A0F0A000"
)
port map (
  I0 => cpi_dbg_data(27),
  I1 => cpi_lddata(27),
  I2 => rst,
  I3 => \GRLFPC20.N_1704\,
  I4 => \GRLFPC20.R.FSR.TEM\(4),
  I5 => \GRLFPC20.N_1338\,
  LO => \GRLFPC20.COMB.V.FSR.TEM_1\(4));
\GRLFPC20.COMB.V.FSR.TEM_1[3]_Z6985\: LUT6_L 
generic map(
  INIT => X"A0C0A0C0A0F0A000"
)
port map (
  I0 => cpi_dbg_data(26),
  I1 => cpi_lddata(26),
  I2 => rst,
  I3 => \GRLFPC20.N_1704\,
  I4 => \GRLFPC20.R.FSR.TEM\(3),
  I5 => \GRLFPC20.N_1338\,
  LO => \GRLFPC20.COMB.V.FSR.TEM_1\(3));
\GRLFPC20.COMB.V.FSR.TEM_1[2]_Z6986\: LUT6_L 
generic map(
  INIT => X"A0C0A0C0A0F0A000"
)
port map (
  I0 => cpi_dbg_data(25),
  I1 => cpi_lddata(25),
  I2 => rst,
  I3 => \GRLFPC20.N_1704\,
  I4 => \GRLFPC20.R.FSR.TEM\(2),
  I5 => \GRLFPC20.N_1338\,
  LO => \GRLFPC20.COMB.V.FSR.TEM_1\(2));
\GRLFPC20.COMB.V.FSR.NONSTD_1_Z6987\: LUT6_L 
generic map(
  INIT => X"A0C0A0C0A0F0A000"
)
port map (
  I0 => cpi_dbg_data(22),
  I1 => cpi_lddata(22),
  I2 => rst,
  I3 => \GRLFPC20.N_1704\,
  I4 => \GRLFPC20.R.FSR.NONSTD\,
  I5 => \GRLFPC20.N_1338\,
  LO => \GRLFPC20.COMB.V.FSR.NONSTD_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[36]_Z6988\: LUT5 
generic map(
  INIT => X"0053FF53"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(23),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(27),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8219\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(36));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[25]\: LUT5 
generic map(
  INIT => X"FACC0ACC"
)
port map (
  I0 => rfo2_data2(29),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(141),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  I4 => \GRLFPC20.FPI.OP2\(32),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7892\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[24]\: LUT5 
generic map(
  INIT => X"FACC0ACC"
)
port map (
  I0 => rfo2_data2(30),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(140),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  I4 => \GRLFPC20.FPI.OP2\(33),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7893\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[21]\: LUT5 
generic map(
  INIT => X"FACA3A0A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(137),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.FPI.OP2\(33),
  I4 => \GRLFPC20.FPI.OP2\(36),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7896\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[18]\: LUT5 
generic map(
  INIT => X"FACA3A0A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(134),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.FPI.OP2\(36),
  I4 => \GRLFPC20.FPI.OP2\(39),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7899\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[16]\: LUT5 
generic map(
  INIT => X"FACA3A0A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(132),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.FPI.OP2\(38),
  I4 => \GRLFPC20.FPI.OP2\(41),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7901\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[15]\: LUT5 
generic map(
  INIT => X"FACA3A0A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(131),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.FPI.OP2\(39),
  I4 => \GRLFPC20.FPI.OP2\(42),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7902\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[14]\: LUT5 
generic map(
  INIT => X"FACA3A0A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(130),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.FPI.OP2\(40),
  I4 => \GRLFPC20.FPI.OP2\(43),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7903\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[9]\: LUT5 
generic map(
  INIT => X"FACA3A0A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(125),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.FPI.OP2\(45),
  I4 => \GRLFPC20.FPI.OP2\(48),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7908\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[8]\: LUT5 
generic map(
  INIT => X"FACA3A0A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(124),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.FPI.OP2\(46),
  I4 => \GRLFPC20.FPI.OP2\(49),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7909\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[7]\: LUT5 
generic map(
  INIT => X"FACA3A0A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(123),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.FPI.OP2\(47),
  I4 => \GRLFPC20.FPI.OP2\(50),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7910\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[3]\: LUT5 
generic map(
  INIT => X"FACA3A0A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(119),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.FPI.OP2\(51),
  I4 => \GRLFPC20.FPI.OP2\(54),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7914\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_14[141]_Z7000\: LUT4_L 
generic map(
  INIT => X"E222"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(143),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_T_3\(0),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_14\(141));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[37]_Z7001\: LUT6 
generic map(
  INIT => X"555500FF33330F0F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(20),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(22),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(26),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(24),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(37));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[35]_Z7002\: LUT6 
generic map(
  INIT => X"555533330F0F00FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(22),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(26),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(24),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(28),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(35));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[33]_Z7003\: LUT5 
generic map(
  INIT => X"530053FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(24),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(28),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8224\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(33));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[31]_Z7004\: LUT5 
generic map(
  INIT => X"0035FF35"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(32),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(28),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8224\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(31));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[29]_Z7005\: LUT5 
generic map(
  INIT => X"350035FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(32),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(28),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8228\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(29));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[22]\: LUT5 
generic map(
  INIT => X"FACA3A0A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(138),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.FPI.OP2\(32),
  I4 => \GRLFPC20.FPI.OP2\(35),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7895\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[20]\: LUT5 
generic map(
  INIT => X"FACA3A0A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(136),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.FPI.OP2\(34),
  I4 => \GRLFPC20.FPI.OP2\(37),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7897\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[19]\: LUT5 
generic map(
  INIT => X"FACA3A0A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(135),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.FPI.OP2\(35),
  I4 => \GRLFPC20.FPI.OP2\(38),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7898\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[17]\: LUT5 
generic map(
  INIT => X"FACA3A0A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(133),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.FPI.OP2\(37),
  I4 => \GRLFPC20.FPI.OP2\(40),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7900\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[13]\: LUT5 
generic map(
  INIT => X"FACA3A0A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(129),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.FPI.OP2\(41),
  I4 => \GRLFPC20.FPI.OP2\(44),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7904\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[11]\: LUT5 
generic map(
  INIT => X"FACA3A0A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(127),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.FPI.OP2\(43),
  I4 => \GRLFPC20.FPI.OP2\(46),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7906\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[10]\: LUT5 
generic map(
  INIT => X"FACA3A0A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(126),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.FPI.OP2\(44),
  I4 => \GRLFPC20.FPI.OP2\(47),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7907\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[6]\: LUT5 
generic map(
  INIT => X"FACA3A0A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(122),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.FPI.OP2\(48),
  I4 => \GRLFPC20.FPI.OP2\(51),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7911\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[5]\: LUT5 
generic map(
  INIT => X"FACA3A0A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(121),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.FPI.OP2\(49),
  I4 => \GRLFPC20.FPI.OP2\(52),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7912\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[4]\: LUT5 
generic map(
  INIT => X"FACA3A0A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(120),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.FPI.OP2\(50),
  I4 => \GRLFPC20.FPI.OP2\(53),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7913\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0[56]_Z7016\: LUT5 
generic map(
  INIT => X"CCCCCAAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(175),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(56));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0[54]_Z7017\: LUT5 
generic map(
  INIT => X"CCCCCAAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(177),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0[38]_Z7018\: LUT5 
generic map(
  INIT => X"CCCCCAAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(193),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(38));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0[37]_Z7019\: LUT5 
generic map(
  INIT => X"CCCCCAAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(194),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(37));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0[36]_Z7020\: LUT5 
generic map(
  INIT => X"CCCCCAAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(195),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(36));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0[33]_Z7021\: LUT5 
generic map(
  INIT => X"CCCCCAAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(198),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(33));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[375]_Z7022\: LUT5_L 
generic map(
  INIT => X"0E0000B0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_2\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(0),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(375));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(259),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(317),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.SI_6\(51));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(274),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(332),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.CIN_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.SI_21\(36));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(272),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(330),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.CIN_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.SI_19\(38));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(271),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(329),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.SI_18\(39));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(269),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(327),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.CIN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.SI_16\(41));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(267),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(325),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.CIN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.SI_14\(43));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(265),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(323),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.SI_12\(45));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(264),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(322),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.CIN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.SI_11\(46));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(263),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(321),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.SI_10\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(262),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(320),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.SI_9\(48));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(261),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(319),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.SI_8\(49));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(290),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(348),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.SI_37\(20));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(289),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(347),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.SI_36\(21));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(287),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(345),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.CIN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.SI_34\(23));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(286),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(344),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.SI_33\(24));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(285),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(343),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.SI_32\(25));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(283),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(341),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.CIN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.SI_30\(27));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(282),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(340),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.CIN_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.SI_29\(28));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(281),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(339),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.CIN_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.SI_28\(29));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(279),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(337),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.SI_26\(31));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(278),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(336),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.SI_25\(32));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(277),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(335),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.CIN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.SI_24\(33));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(276),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(334),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.SI_23\(34));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(298),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(356),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.SI_45\(12));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43.Z_AXBXC0\: LUT4 
generic map(
  INIT => X"2DD2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(355),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(18),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.SI_44\(13));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(296),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(354),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.SI_43\(14));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39.Z_AXBXC0\: LUT4 
generic map(
  INIT => X"2DD2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(351),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(22),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.CIN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.SI_40\(17));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"0F660066F099FF99"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(292),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(350),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.SI_39\(18));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(304),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(362),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.CIN_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.SI_51\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(303),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(361),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.SI_50\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(300),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(358),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.SI_47\(10));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(309),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(367),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.SI_56\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53.Z_AXBXC0\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(307),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(365),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.SI_54\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNICFTG1[229]\: LUT6 
generic map(
  INIT => X"CC33CC33CA35AC53"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(229),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => N_6674);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIADTG1[228]\: LUT6 
generic map(
  INIT => X"CC33CC33CA35AC53"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(228),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => N_6682);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI8BTG1[227]\: LUT6 
generic map(
  INIT => X"CC33CC33CA35AC53"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(227),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => N_6690);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[374]_Z7059\: LUT5_L 
generic map(
  INIT => X"01FFFF40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_2\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(0),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(374));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT_Z7060\: LUT5 
generic map(
  INIT => X"F4000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CONDMUXMULXFF.UN5_NOTSQRTLFTCC\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_WQSTSETS\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6[53]_Z7061\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFFF20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2229_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_906\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9972_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10304\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(53),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_0\(53),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(53));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_1[48]_Z7062\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF0040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10146\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12021_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_795\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10164\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(48),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_1\(48));
\GRLFPC20.COMB.V.I.RES_1[50]_Z7063\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(50),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(53),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.FRAC\(53),
  LO => \GRLFPC20.COMB.V.I.RES_1\(50));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.OPREXCSHFT.UN3_OPREXC_Z7064\: LUT5 
generic map(
  INIT => X"FFFE0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(248),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(249),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(247),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1_3\(6),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\(4),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.OPREXCSHFT.UN3_OPREXC\);
\GRLFPC20.COMB.V.E.STDATA_1[20]_Z7065\: LUT6_L 
generic map(
  INIT => X"E400E4FFE400E400"
)
port map (
  I0 => \GRLFPC20.COMB.V.E.STDATA2\,
  I1 => \GRLFPC20.R.I.INST\(20),
  I2 => \GRLFPC20.R.I.PC\(20),
  I3 => \GRLFPC20.R.A.AFQ\,
  I4 => \GRLFPC20.R.A.AFSR\,
  I5 => \GRLFPC20.FPI.OP1\(52),
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(20));
\GRLFPC20.COMB.V.I.RES_1[55]_Z7066\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(55),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(58),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.EXP\(3),
  LO => \GRLFPC20.COMB.V.I.RES_1\(55));
\GRLFPC20.COMB.V.E.STDATA_1[29]_Z7067\: LUT6_L 
generic map(
  INIT => X"D800D8FFD800D800"
)
port map (
  I0 => \GRLFPC20.COMB.V.E.STDATA2\,
  I1 => \GRLFPC20.R.I.PC\(29),
  I2 => \GRLFPC20.R.I.INST\(29),
  I3 => \GRLFPC20.R.A.AFQ\,
  I4 => \GRLFPC20.R.A.AFSR\,
  I5 => \GRLFPC20.FPI.OP1\(61),
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(29));
\GRLFPC20.COMB.V.I.RES_1[57]_Z7068\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(57),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(60),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.EXP\(5),
  LO => \GRLFPC20.COMB.V.I.RES_1\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL[67]_Z7069\: LUT5 
generic map(
  INIT => X"00020202"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(47),
  I1 => \GRLFPC20.FPI.LDOP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(12),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS\,
  I4 => N_3882,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67));
\GRLFPC20.COMB.V.I.RES_1[31]_Z7070\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(31),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(34),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.FRAC\(34),
  LO => \GRLFPC20.COMB.V.I.RES_1\(31));
\GRLFPC20.WRADDR_1[2]\: LUT6 
generic map(
  INIT => X"AAAAAAAACCCFCCC0"
)
port map (
  I0 => cpi_dbg_addr(2),
  I1 => cpi_x_inst(27),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.UN1_R.I.V\,
  I4 => \GRLFPC20.R.I.INST\(27),
  I5 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => RFI2_WRADDR_25);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1[34]_Z7072\: LUT4 
generic map(
  INIT => X"0028"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\(34));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1[35]_Z7073\: LUT4 
generic map(
  INIT => X"0028"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\(35));
\GRLFPC20.WRADDR_1[4]\: LUT6 
generic map(
  INIT => X"AAAAAAAACCCFCCC0"
)
port map (
  I0 => cpi_dbg_addr(4),
  I1 => cpi_x_inst(29),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.UN1_R.I.V\,
  I4 => \GRLFPC20.R.I.INST\(29),
  I5 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => RFI2_WRADDR_27);
\GRLFPC20.COMB.V.E.STDATA_1[17]_Z7075\: LUT6_L 
generic map(
  INIT => X"E4FFE4FFE4FFE400"
)
port map (
  I0 => \GRLFPC20.COMB.V.E.STDATA2\,
  I1 => \GRLFPC20.R.I.INST\(17),
  I2 => \GRLFPC20.R.I.PC\(17),
  I3 => \GRLFPC20.R.A.AFQ\,
  I4 => \GRLFPC20.R.A.AFSR\,
  I5 => \GRLFPC20.FPI.OP1\(49),
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(17));
\GRLFPC20.COMB.V.E.STDATA_1[21]_Z7076\: LUT6_L 
generic map(
  INIT => X"E400E4FFE400E400"
)
port map (
  I0 => \GRLFPC20.COMB.V.E.STDATA2\,
  I1 => \GRLFPC20.R.I.INST\(21),
  I2 => \GRLFPC20.R.I.PC\(21),
  I3 => \GRLFPC20.R.A.AFQ\,
  I4 => \GRLFPC20.R.A.AFSR\,
  I5 => \GRLFPC20.FPI.OP1\(53),
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(21));
\GRLFPC20.WRADDR_1[1]\: LUT6 
generic map(
  INIT => X"AAAAAAAACCCFCCC0"
)
port map (
  I0 => cpi_dbg_addr(1),
  I1 => cpi_x_inst(26),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.UN1_R.I.V\,
  I4 => \GRLFPC20.R.I.INST\(26),
  I5 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => RFI2_WRADDR_24);
\GRLFPC20.WRADDR_1[3]\: LUT6 
generic map(
  INIT => X"AAAAAAAACCCFCCC0"
)
port map (
  I0 => cpi_dbg_addr(3),
  I1 => cpi_x_inst(28),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.COMB.UN1_R.I.V\,
  I4 => \GRLFPC20.R.I.INST\(28),
  I5 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => RFI2_WRADDR_26);
\GRLFPC20.COMB.V.I.RES_1[29]_Z7079\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(29),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(32),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.FRAC\(32),
  LO => \GRLFPC20.COMB.V.I.RES_1\(29));
\GRLFPC20.COMB.V.I.RES_1[30]_Z7080\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(30),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(33),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.FRAC\(33),
  LO => \GRLFPC20.COMB.V.I.RES_1\(30));
\GRLFPC20.COMB.V.I.RES_1[32]_Z7081\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(32),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(35),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.FRAC\(35),
  LO => \GRLFPC20.COMB.V.I.RES_1\(32));
\GRLFPC20.COMB.V.I.RES_1[33]_Z7082\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(33),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(36),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.FRAC\(36),
  LO => \GRLFPC20.COMB.V.I.RES_1\(33));
\GRLFPC20.COMB.V.I.RES_1[34]_Z7083\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(34),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(37),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.FRAC\(37),
  LO => \GRLFPC20.COMB.V.I.RES_1\(34));
\GRLFPC20.COMB.V.I.RES_1[35]_Z7084\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(35),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(38),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.FRAC\(38),
  LO => \GRLFPC20.COMB.V.I.RES_1\(35));
\GRLFPC20.COMB.V.I.RES_1[36]_Z7085\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(36),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(39),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.FRAC\(39),
  LO => \GRLFPC20.COMB.V.I.RES_1\(36));
\GRLFPC20.COMB.V.I.RES_1[37]_Z7086\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(37),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(40),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.FRAC\(40),
  LO => \GRLFPC20.COMB.V.I.RES_1\(37));
\GRLFPC20.COMB.V.I.RES_1[38]_Z7087\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(38),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(41),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.FRAC\(41),
  LO => \GRLFPC20.COMB.V.I.RES_1\(38));
\GRLFPC20.COMB.V.I.RES_1[39]_Z7088\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(39),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(42),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.FRAC\(42),
  LO => \GRLFPC20.COMB.V.I.RES_1\(39));
\GRLFPC20.COMB.V.I.RES_1[40]_Z7089\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(40),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(43),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.FRAC\(43),
  LO => \GRLFPC20.COMB.V.I.RES_1\(40));
\GRLFPC20.COMB.V.I.RES_1[41]_Z7090\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(41),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(44),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.FRAC\(44),
  LO => \GRLFPC20.COMB.V.I.RES_1\(41));
\GRLFPC20.COMB.V.I.RES_1[42]_Z7091\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(42),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(45),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.FRAC\(45),
  LO => \GRLFPC20.COMB.V.I.RES_1\(42));
\GRLFPC20.COMB.V.I.RES_1[43]_Z7092\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(43),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(46),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.FRAC\(46),
  LO => \GRLFPC20.COMB.V.I.RES_1\(43));
\GRLFPC20.COMB.V.I.RES_1[44]_Z7093\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(44),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(47),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.FRAC\(47),
  LO => \GRLFPC20.COMB.V.I.RES_1\(44));
\GRLFPC20.COMB.V.I.RES_1[45]_Z7094\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(45),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(48),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.FRAC\(48),
  LO => \GRLFPC20.COMB.V.I.RES_1\(45));
\GRLFPC20.COMB.V.I.RES_1[46]_Z7095\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(46),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(49),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.FRAC\(49),
  LO => \GRLFPC20.COMB.V.I.RES_1\(46));
\GRLFPC20.COMB.V.I.RES_1[47]_Z7096\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(47),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(50),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.FRAC\(50),
  LO => \GRLFPC20.COMB.V.I.RES_1\(47));
\GRLFPC20.COMB.V.I.RES_1[48]_Z7097\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(48),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(51),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.FRAC\(51),
  LO => \GRLFPC20.COMB.V.I.RES_1\(48));
\GRLFPC20.COMB.V.I.RES_1[49]_Z7098\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(49),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(52),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.FRAC\(52),
  LO => \GRLFPC20.COMB.V.I.RES_1\(49));
\GRLFPC20.COMB.V.I.RES_1[51]_Z7099\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(51),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(54),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.FRAC\(54),
  LO => \GRLFPC20.COMB.V.I.RES_1\(51));
\GRLFPC20.COMB.V.I.RES_1[52]_Z7100\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(52),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(55),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.EXP\(0),
  LO => \GRLFPC20.COMB.V.I.RES_1\(52));
\GRLFPC20.COMB.V.I.RES_1[53]_Z7101\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(53),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(56),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.EXP\(1),
  LO => \GRLFPC20.COMB.V.I.RES_1\(53));
\GRLFPC20.COMB.V.I.RES_1[54]_Z7102\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(54),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(57),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.EXP\(2),
  LO => \GRLFPC20.COMB.V.I.RES_1\(54));
\GRLFPC20.COMB.V.I.RES_1[56]_Z7103\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(56),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(59),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.EXP\(4),
  LO => \GRLFPC20.COMB.V.I.RES_1\(56));
\GRLFPC20.COMB.V.I.RES_1[58]_Z7104\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(58),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(61),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.EXP\(6),
  LO => \GRLFPC20.COMB.V.I.RES_1\(58));
\GRLFPC20.COMB.V.I.RES_1[59]_Z7105\: LUT5_L 
generic map(
  INIT => X"F3E2C0E2"
)
port map (
  I0 => \GRLFPC20.R.I.RES\(59),
  I1 => \GRLFPC20.N_1858\,
  I2 => \GRLFPC20.FPI.OP2\(62),
  I3 => \GRLFPC20.N_2102\,
  I4 => \GRLFPC20.FPO.EXP\(7),
  LO => \GRLFPC20.COMB.V.I.RES_1\(59));
\GRLFPC20.COMB.V.E.STDATA_1[12]_Z7106\: LUT6_L 
generic map(
  INIT => X"E400E4FFE400E400"
)
port map (
  I0 => \GRLFPC20.COMB.V.E.STDATA2\,
  I1 => \GRLFPC20.R.I.INST\(12),
  I2 => \GRLFPC20.R.I.PC\(12),
  I3 => \GRLFPC20.R.A.AFQ\,
  I4 => \GRLFPC20.R.A.AFSR\,
  I5 => \GRLFPC20.FPI.OP1\(44),
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(12));
\GRLFPC20.COMB.V.E.STDATA_1[18]_Z7107\: LUT6_L 
generic map(
  INIT => X"E4FFE4FFE4FFE400"
)
port map (
  I0 => \GRLFPC20.COMB.V.E.STDATA2\,
  I1 => \GRLFPC20.R.I.INST\(18),
  I2 => \GRLFPC20.R.I.PC\(18),
  I3 => \GRLFPC20.R.A.AFQ\,
  I4 => \GRLFPC20.R.A.AFSR\,
  I5 => \GRLFPC20.FPI.OP1\(50),
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(18));
\GRLFPC20.COMB.V.E.STDATA_1[19]_Z7108\: LUT6_L 
generic map(
  INIT => X"D800D8FFD800D800"
)
port map (
  I0 => \GRLFPC20.COMB.V.E.STDATA2\,
  I1 => \GRLFPC20.R.I.PC\(19),
  I2 => \GRLFPC20.R.I.INST\(19),
  I3 => \GRLFPC20.R.A.AFQ\,
  I4 => \GRLFPC20.R.A.AFSR\,
  I5 => \GRLFPC20.FPI.OP1\(51),
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(19));
\GRLFPC20.COMB.V.E.STDATA_1[28]_Z7109\: LUT6_L 
generic map(
  INIT => X"D800D8FFD800D800"
)
port map (
  I0 => \GRLFPC20.COMB.V.E.STDATA2\,
  I1 => \GRLFPC20.R.I.PC\(28),
  I2 => \GRLFPC20.R.I.INST\(28),
  I3 => \GRLFPC20.R.A.AFQ\,
  I4 => \GRLFPC20.R.A.AFSR\,
  I5 => \GRLFPC20.FPI.OP1\(60),
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(28));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1[33]_Z7110\: LUT4 
generic map(
  INIT => X"0028"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\(33));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1[36]_Z7111\: LUT4 
generic map(
  INIT => X"0028"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\(36));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1[37]_Z7112\: LUT4 
generic map(
  INIT => X"0028"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\(37));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1[38]_Z7113\: LUT4 
generic map(
  INIT => X"0028"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\(38));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_DIVMULTV[0]_Z7114\: LUT4_L 
generic map(
  INIT => X"4002"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(3),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(2),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(0),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_DIVMULTV\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1[54]_Z7115\: LUT4 
generic map(
  INIT => X"0028"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[2]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF7350"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1006_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2730\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2565\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2502\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[14]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF20FF2020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_742\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2600\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2730\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0\(14),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(14));
\GRLFPC20.COMB.SEQERR.UN11_OP\: LUT6 
generic map(
  INIT => X"0000000B00000000"
)
port map (
  I0 => cpi_d_inst(19),
  I1 => cpi_d_inst(20),
  I2 => cpi_d_inst(21),
  I3 => cpi_d_inst(22),
  I4 => cpi_d_inst(23),
  I5 => cpi_d_inst(24),
  O => \GRLFPC20.N_1142\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.ENTRYPOINT_Z7119\: LUT6 
generic map(
  INIT => X"00000000000051F3"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9913_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_9_0\(47),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN1_S_14\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN3_S_SQRT_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN10_S_MOV\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(45),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.ENTRYPOINT\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[43]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFEAC0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2584\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10246_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2608\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2758\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2216\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1653\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(43));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5[61]_Z7121\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF8000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9549_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9994_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10869\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10888_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_0\(61),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2\(61),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5\(61));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2[23]_Z7122\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFF8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2762\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(23),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2400\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2403\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1039\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2\(23));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1[26]_Z7123\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF80B0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2645\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9558_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2583\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_717\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2380\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_1\(26),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1\(26));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0[29]_Z7124\: LUT6 
generic map(
  INIT => X"FFFFFFFFF111F000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_741\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1335\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_777\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1169\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_866\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(29));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2[3]_Z7125\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10592_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2600\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2563\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2129\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6[36]_Z7126\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFFFF2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9922_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12195\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10022\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10024\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_0\(36),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_1\(36),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(36));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_0[27]_Z7127\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9968_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9790_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10790\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_783\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9794\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0\(27),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_0\(27));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7[27]_Z7128\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF3222"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9800_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10410\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10943\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9801\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0\(27),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7\(27));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4[13]_Z7129\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFF10000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_125\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9389_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_10_1\(61),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9671_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10943\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_1\(13),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4\(13));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_0[4]_Z7130\: LUT6 
generic map(
  INIT => X"FFFFFFFF2F222222"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_7_0\(4),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_85\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9911_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9506_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10246_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(4),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_0\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1[4]_Z7131\: LUT5 
generic map(
  INIT => X"FFFFFFF8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_0\(11),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2583\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2831\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2335\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_0\(4),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1[50]_Z7132\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF8F88"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_6081_A2_6_0\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2701\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10410\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1282\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2156\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1654\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1\(50));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_0[7]_Z7133\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1553_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_749\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_291_I\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2219\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(7),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_0\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1[7]_Z7134\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFFF40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_783\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2584\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10943\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2224\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2512\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_0\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6[48]_Z7135\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF04"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9887_I\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10161_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_795\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10166\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10167\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3\(48),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(48));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8[55]_Z7136\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFFF08"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9700_I\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10479\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_289\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10446\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3\(55),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(55),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8\(55));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9[55]_Z7137\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF08"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2635\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9604_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10025_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10458\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10460\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5\(55),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9\(55));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_0[59]_Z7138\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_767_I\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9915_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10752_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_1\(59),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0\(59),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(59),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_0\(59));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0[32]_Z7139\: LUT6_L 
generic map(
  INIT => X"083B080800000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1561\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9508_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9828\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9338_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_6_1\(32),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0\(32));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1[12]_Z7140\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFEAC0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_0\(4),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_134_I\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2842\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1711\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1648\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1\(12));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_7_0[11]_Z7141\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFF2F0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10640\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_741\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9328\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9604_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9314\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2\(11),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_7_0\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_1_1[11]_Z7142\: LUT4_L 
generic map(
  INIT => X"FFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12250\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_5_0\(11),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9338\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_6\(11),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_1_1\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_6_0[31]_Z7143\: LUT6 
generic map(
  INIT => X"FFFFFFFFA0A0ECA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9428\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9390_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9404_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10888_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9785_1_I_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_1_0\(31),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_6_0\(31));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_7_0[31]_Z7144\: LUT6 
generic map(
  INIT => X"FFFFFFFF00A0CCEC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9600_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1149\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1175\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_720\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_765\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_3_0\(31),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_7_0\(31));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_0_1[31]_Z7145\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF10"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9629\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_906\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9916_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_4_1\(31),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9409\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_5\(31),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_0_1\(31));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7[6]_Z7146\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF08"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9505_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9738_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2167\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_1\(6),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3\(6),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_0[17]_Z7147\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFFF80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10592_I\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9558_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2584\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2445\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_979\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_978\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_0\(17));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4[19]_Z7148\: LUT6 
generic map(
  INIT => X"FFFFDCCC50005000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_796\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_8_1\(19),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9670_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9604_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_3_2\(19),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6[19]_Z7149\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF00D0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_766\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9604_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9394_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_720\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9652\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_1\(19),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8[19]_Z7150\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF0080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9657_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1132_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_314_I\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3\(19),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0\(19),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8[33]_Z7151\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9906_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10888_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9666_1_I_0\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9971\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_1\(33),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4\(33),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8\(33));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6[58]_Z7152\: LUT6 
generic map(
  INIT => X"FFFFFFFF75553000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_907\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9994_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1149\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10631_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10694_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(58),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(58));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7_1[58]_Z7153\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFCECC0A00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1149\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10661\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_409\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_995_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10243_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(58),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7_1\(58));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8_2[58]_Z7154\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10670_I\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9973_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9671_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0\(58),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_981\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9453\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8_2\(58));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9[58]_Z7155\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF88F8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10693_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_291_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1232\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12131\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4\(58),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_1\(58),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9\(58));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9[54]_Z7156\: LUT6 
generic map(
  INIT => X"FFFFFFFFECCCA000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2669\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_10_1\(61),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_795\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9453_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10943\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9_0\(54),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0[54]_Z7157\: LUT6 
generic map(
  INIT => X"FFFFFFFFFF040404"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10343_I\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9797_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_795\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9604_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2591\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(54),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_5[56]_Z7158\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFF8FFF0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_732\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_0\(56),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1009\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1002_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10531\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_5\(56));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_0[51]_Z7159\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFAAEA00C0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_2_A2_0_A2_0\(51),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9700_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10891_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_328\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2584\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(51),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_0\(51));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_4_1[51]_Z7160\: LUT6 
generic map(
  INIT => X"FFFFFFFFCE0ACC00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_0_A2_0_A2_0\(51),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10584_I\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2600\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1282\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_0\(51),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_4_1\(51));
\GRLFPC20.R.I.RDD_RNO\: LUT6_L 
generic map(
  INIT => X"2200AA002020A0A0"
)
port map (
  I0 => rst,
  I1 => \GRLFPC20.R.A.MOV\,
  I2 => \GRLFPC20.R.I.RDD\,
  I3 => \GRLFPC20.R.X.RDD\,
  I4 => \GRLFPC20.N_2931_1\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  LO => \GRLFPC20.N_3022_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_1_O2[37]\: LUT6 
generic map(
  INIT => X"FFFFFFFF0F0F0400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_732\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_291_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9666_1_I_0\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1157\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2255\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_782\);
\GRLFPC20.RS1D_CNST.M6\: LUT6 
generic map(
  INIT => X"0810080008000800"
)
port map (
  I0 => cpi_d_inst(19),
  I1 => cpi_d_inst(20),
  I2 => cpi_d_inst(23),
  I3 => cpi_d_inst(30),
  I4 => \GRLFPC20.N_3116\,
  I5 => \GRLFPC20.N_3128\,
  O => \GRLFPC20.RS1D_CNST.N_7\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_11[75]\: LUT5 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(49),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(51),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8807\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8810\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8814\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8815\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_WQSTSETS[0]_Z7165\: LUT6 
generic map(
  INIT => X"0004000433370004"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_I_I_A2_0_O2_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_SM12\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN11_WQSTSETS_0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_WQSTSETS\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI0HPS3[59]\: LUT6 
generic map(
  INIT => X"C33CA55AF0F0F0F0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_AXB0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_I_20\: LUT6_L 
generic map(
  INIT => X"E01F20DF1FE0DF20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(236),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1137\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(8),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12036\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_RNINJCT3[57]\: LUT6 
generic map(
  INIT => X"C33C699633CC33CC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(57),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIAML61[311]\: LUT6 
generic map(
  INIT => X"F099FF990F660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(311),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(369),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SALSBS_1\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0[61]_Z7170\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF0002"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9555_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10824_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_831\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10869\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10892\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10884\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(61));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1[34]_Z7171\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFFF80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9739_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12021_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9972_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9971\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9969\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9968\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(34));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_RNIH63D1\: LUT6 
generic map(
  INIT => X"AC00FFFF53FF0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN16_NOTPROP_2336_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19[70]_Z7173\: LUT6 
generic map(
  INIT => X"FF00F0F0CCCCAAAA"
)
port map (
  I0 => rfo1_data1(10),
  I1 => rfo1_data1(13),
  I2 => rfo2_data1(10),
  I3 => rfo2_data1(13),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I5 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(70));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19[77]_Z7174\: LUT5 
generic map(
  INIT => X"FC0CFA0A"
)
port map (
  I0 => rfo1_data1(3),
  I1 => rfo2_data1(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.OP1\(38),
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(77));
\GRLFPC20.COMB.V.E.STDATA_1_1[23]\: LUT5_L 
generic map(
  INIT => X"F0CCF0AA"
)
port map (
  I0 => rfo1_data1(23),
  I1 => rfo2_data1(23),
  I2 => \GRLFPC20.R.FSR.TEM\(0),
  I3 => \GRLFPC20.R.A.AFSR\,
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  LO => \GRLFPC20.N_2395\);
\GRLFPC20.COMB.RS1_1_1[0]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => cpi_d_inst(25),
  I1 => \GRLFPC20.RS1V_0_SQMUXA\,
  O => \GRLFPC20.N_2512\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[43]\: LUT6 
generic map(
  INIT => X"00FF0F0F33335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8212\);
\GRLFPC20.COMB.V.E.STDATA_1_1[25]\: LUT5_L 
generic map(
  INIT => X"F0CCF0AA"
)
port map (
  I0 => rfo1_data1(25),
  I1 => rfo2_data1(25),
  I2 => \GRLFPC20.R.FSR.TEM\(2),
  I3 => \GRLFPC20.R.A.AFSR\,
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  LO => \GRLFPC20.N_2397\);
\GRLFPC20.COMB.V.E.STDATA_1_1[16]\: LUT5_L 
generic map(
  INIT => X"F0CCF0AA"
)
port map (
  I0 => rfo1_data1(16),
  I1 => rfo2_data1(16),
  I2 => \GRLFPC20.R.FSR.FTT\(2),
  I3 => \GRLFPC20.R.A.AFSR\,
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  LO => \GRLFPC20.N_2388\);
\GRLFPC20.COMB.V.E.STDATA_1_1[13]\: LUT6_L 
generic map(
  INIT => X"00F0CCCC00F0AAAA"
)
port map (
  I0 => rfo1_data1(13),
  I1 => rfo2_data1(13),
  I2 => \GRLFPC20.R.STATE\(1),
  I3 => \GRLFPC20.R.STATE\(0),
  I4 => \GRLFPC20.R.A.AFSR\,
  I5 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  LO => \GRLFPC20.N_2385\);
\GRLFPC20.COMB.V.FSR.TEM_1[0]_Z7181\: LUT6_L 
generic map(
  INIT => X"A0C0A0C0A0F0A000"
)
port map (
  I0 => cpi_dbg_data(23),
  I1 => cpi_lddata(23),
  I2 => rst,
  I3 => \GRLFPC20.N_1704\,
  I4 => \GRLFPC20.R.FSR.TEM\(0),
  I5 => \GRLFPC20.N_1338\,
  LO => \GRLFPC20.COMB.V.FSR.TEM_1\(0));
\GRLFPC20.COMB.V.FSR.TEM_1[1]_Z7182\: LUT6_L 
generic map(
  INIT => X"A0C0A0C0A0F0A000"
)
port map (
  I0 => cpi_dbg_data(24),
  I1 => cpi_lddata(24),
  I2 => rst,
  I3 => \GRLFPC20.N_1704\,
  I4 => \GRLFPC20.R.FSR.TEM\(1),
  I5 => \GRLFPC20.N_1338\,
  LO => \GRLFPC20.COMB.V.FSR.TEM_1\(1));
\GRLFPC20.COMB.V.FSR.RD_1[1]_Z7183\: LUT6_L 
generic map(
  INIT => X"A0C0A0C0A0F0A000"
)
port map (
  I0 => cpi_dbg_data(31),
  I1 => cpi_lddata(31),
  I2 => rst,
  I3 => \GRLFPC20.N_1704\,
  I4 => \GRLFPC20.R.FSR.RD\(1),
  I5 => \GRLFPC20.N_1338\,
  LO => \GRLFPC20.COMB.V.FSR.RD_1\(1));
\GRLFPC20.COMB.V.FSR.RD_1[0]_Z7184\: LUT6_L 
generic map(
  INIT => X"A0C0A0C0A0F0A000"
)
port map (
  I0 => cpi_dbg_data(30),
  I1 => cpi_lddata(30),
  I2 => rst,
  I3 => \GRLFPC20.N_1704\,
  I4 => \GRLFPC20.R.FSR.RD\(0),
  I5 => \GRLFPC20.N_1338\,
  LO => \GRLFPC20.COMB.V.FSR.RD_1\(0));
\GRLFPC20.WRDATA[63]\: LUT5 
generic map(
  INIT => X"AAAACFC0"
)
port map (
  I0 => cpi_dbg_data(31),
  I1 => cpi_lddata(31),
  I2 => \GRLFPC20.N_1562\,
  I3 => \GRLFPC20.R.I.RES\(63),
  I4 => \GRLFPC20.WRADDR_0_SQMUXA\,
  O => rfi1_wrdata(31));
\GRLFPC20.COMB.LOCKGEN.UN7_DEPCHECK\: LUT6 
generic map(
  INIT => X"EEEEEEEEEEEEEEE0"
)
port map (
  I0 => \GRLFPC20.COMB.FPDECODE.ST\,
  I1 => \GRLFPC20.N_1583\,
  I2 => \GRLFPC20.R.A.LD\,
  I3 => \GRLFPC20.R.E.LD\,
  I4 => \GRLFPC20.R.M.LD\,
  I5 => \GRLFPC20.R.X.LD\,
  O => \GRLFPC20.N_1597\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[25]\: LUT6 
generic map(
  INIT => X"00FF33330F0F5555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8230\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[37]\: LUT6 
generic map(
  INIT => X"0F0F3333555500FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8218\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[18]\: LUT6 
generic map(
  INIT => X"0F0F00FF55553333"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8237\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[20]\: LUT6 
generic map(
  INIT => X"00FF33330F0F5555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8235\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[24]\: LUT6 
generic map(
  INIT => X"00FF0F0F55553333"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8231\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[40]\: LUT6 
generic map(
  INIT => X"333300FF0F0F5555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8215\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[44]\: LUT6 
generic map(
  INIT => X"00FF55550F0F3333"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8211\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[17]\: LUT6 
generic map(
  INIT => X"00FF0F0F55553333"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8238\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[21]\: LUT6 
generic map(
  INIT => X"0F0F00FF33335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8234\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[57]\: LUT6 
generic map(
  INIT => X"00FF0F0F33335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8198\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[56]\: LUT6 
generic map(
  INIT => X"00FF0F0F55553333"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8199\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[55]\: LUT6 
generic map(
  INIT => X"00FF0F0F33335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8200\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[54]\: LUT6 
generic map(
  INIT => X"00FF0F0F33335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8201\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[53]\: LUT6 
generic map(
  INIT => X"00FF0F0F33335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8202\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[52]\: LUT6 
generic map(
  INIT => X"00FF33330F0F5555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8203\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[51]\: LUT6 
generic map(
  INIT => X"00FF0F0F33335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8204\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[50]\: LUT6 
generic map(
  INIT => X"00FF0F0F55553333"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8205\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[49]\: LUT6 
generic map(
  INIT => X"00FF0F0F55553333"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8206\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[48]\: LUT6 
generic map(
  INIT => X"0F0F00FF55553333"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8207\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[46]\: LUT6 
generic map(
  INIT => X"00FF33330F0F5555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8209\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[45]\: LUT6 
generic map(
  INIT => X"00FF33330F0F5555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8210\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[41]\: LUT6 
generic map(
  INIT => X"0F0F00FF33335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8214\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[22]\: LUT6 
generic map(
  INIT => X"00FF33330F0F5555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8233\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[19]\: LUT6 
generic map(
  INIT => X"00FF33330F0F5555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8236\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[23]\: LUT6 
generic map(
  INIT => X"0F0F00FF55553333"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8232\);
\GRLFPC20.COMB.V.E.STDATA_1_1[31]\: LUT5_L 
generic map(
  INIT => X"F0CCF0AA"
)
port map (
  I0 => rfo1_data1(31),
  I1 => rfo2_data1(31),
  I2 => \GRLFPC20.R.FSR.RD\(1),
  I3 => \GRLFPC20.R.A.AFSR\,
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  LO => \GRLFPC20.N_2403\);
\GRLFPC20.COMB.V.E.STDATA_1_1[14]\: LUT5_L 
generic map(
  INIT => X"F0CCF0AA"
)
port map (
  I0 => rfo1_data1(14),
  I1 => rfo2_data1(14),
  I2 => \GRLFPC20.R.FSR.FTT\(0),
  I3 => \GRLFPC20.R.A.AFSR\,
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  LO => \GRLFPC20.N_2386\);
\GRLFPC20.COMB.V.E.STDATA_1_1[2]\: LUT5_L 
generic map(
  INIT => X"F0CCF0AA"
)
port map (
  I0 => rfo1_data1(2),
  I1 => rfo2_data1(2),
  I2 => \GRLFPC20.R.FSR.CEXC\(2),
  I3 => \GRLFPC20.R.A.AFSR\,
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  LO => \GRLFPC20.N_2374\);
\GRLFPC20.COMB.V.E.STDATA_1_1[3]\: LUT5_L 
generic map(
  INIT => X"F0CCF0AA"
)
port map (
  I0 => rfo1_data1(3),
  I1 => rfo2_data1(3),
  I2 => \GRLFPC20.R.FSR.CEXC\(3),
  I3 => \GRLFPC20.R.A.AFSR\,
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  LO => \GRLFPC20.N_2375\);
\GRLFPC20.COMB.V.E.STDATA_1_1[5]\: LUT5_L 
generic map(
  INIT => X"F0CCF0AA"
)
port map (
  I0 => rfo1_data1(5),
  I1 => rfo2_data1(5),
  I2 => \GRLFPC20.R.FSR.AEXC\(0),
  I3 => \GRLFPC20.R.A.AFSR\,
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  LO => \GRLFPC20.N_2377\);
\GRLFPC20.COMB.V.E.STDATA_1_1[7]\: LUT5_L 
generic map(
  INIT => X"F0CCF0AA"
)
port map (
  I0 => rfo1_data1(7),
  I1 => rfo2_data1(7),
  I2 => \GRLFPC20.R.FSR.AEXC\(2),
  I3 => \GRLFPC20.R.A.AFSR\,
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  LO => \GRLFPC20.N_2379\);
\GRLFPC20.COMB.V.E.STDATA_1_1[9]\: LUT5_L 
generic map(
  INIT => X"F0CCF0AA"
)
port map (
  I0 => rfo1_data1(9),
  I1 => rfo2_data1(9),
  I2 => \GRLFPC20.R.FSR.AEXC\(4),
  I3 => \GRLFPC20.R.A.AFSR\,
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  LO => \GRLFPC20.N_2381\);
\GRLFPC20.COMB.V.E.STDATA_1_1[10]\: LUT5_L 
generic map(
  INIT => X"F0CCF0AA"
)
port map (
  I0 => rfo1_data1(10),
  I1 => rfo2_data1(10),
  I2 => NN_1,
  I3 => \GRLFPC20.R.A.AFSR\,
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  LO => \GRLFPC20.N_2382\);
\GRLFPC20.COMB.V.E.STDATA_1_1[11]\: LUT5_L 
generic map(
  INIT => X"F0CCF0AA"
)
port map (
  I0 => rfo1_data1(11),
  I1 => rfo2_data1(11),
  I2 => CPO_CC_3,
  I3 => \GRLFPC20.R.A.AFSR\,
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  LO => \GRLFPC20.N_2383\);
\GRLFPC20.COMB.V.E.STDATA_1_1[24]\: LUT5_L 
generic map(
  INIT => X"F0CCF0AA"
)
port map (
  I0 => rfo1_data1(24),
  I1 => rfo2_data1(24),
  I2 => \GRLFPC20.R.FSR.TEM\(1),
  I3 => \GRLFPC20.R.A.AFSR\,
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  LO => \GRLFPC20.N_2396\);
\GRLFPC20.COMB.V.E.STDATA_1_1[26]\: LUT5_L 
generic map(
  INIT => X"F0CCF0AA"
)
port map (
  I0 => rfo1_data1(26),
  I1 => rfo2_data1(26),
  I2 => \GRLFPC20.R.FSR.TEM\(3),
  I3 => \GRLFPC20.R.A.AFSR\,
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  LO => \GRLFPC20.N_2398\);
\GRLFPC20.COMB.V.E.STDATA_1_1[27]\: LUT5_L 
generic map(
  INIT => X"F0CCF0AA"
)
port map (
  I0 => rfo1_data1(27),
  I1 => rfo2_data1(27),
  I2 => \GRLFPC20.R.FSR.TEM\(4),
  I3 => \GRLFPC20.R.A.AFSR\,
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  LO => \GRLFPC20.N_2399\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19[80]_Z7224\: LUT5 
generic map(
  INIT => X"CFC0AFA0"
)
port map (
  I0 => rfo1_data1(3),
  I1 => rfo2_data1(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.OP1\(32),
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(80));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19[78]_Z7225\: LUT6 
generic map(
  INIT => X"FF00F0F0CCCCAAAA"
)
port map (
  I0 => rfo1_data1(2),
  I1 => rfo1_data1(5),
  I2 => rfo2_data1(2),
  I3 => rfo2_data1(5),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I5 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(78));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19[74]_Z7226\: LUT5 
generic map(
  INIT => X"CFC0AFA0"
)
port map (
  I0 => rfo1_data1(9),
  I1 => rfo2_data1(9),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.OP1\(38),
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(74));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19[67]_Z7227\: LUT6 
generic map(
  INIT => X"FF00F0F0CCCCAAAA"
)
port map (
  I0 => rfo1_data1(13),
  I1 => rfo1_data1(16),
  I2 => rfo2_data1(13),
  I3 => rfo2_data1(16),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I5 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(67));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[47]\: LUT6 
generic map(
  INIT => X"00FF0F0F33335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8208\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[42]\: LUT6 
generic map(
  INIT => X"0F0F00FF33335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8213\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[39]\: LUT6 
generic map(
  INIT => X"00FF0F0F33335555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8216\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[36]\: LUT6 
generic map(
  INIT => X"0F0F3333555500FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8219\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[32]\: LUT6 
generic map(
  INIT => X"3333555500FF0F0F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8223\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[28]\: LUT6 
generic map(
  INIT => X"333300FF0F0F5555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8227\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15[3]\: LUT6 
generic map(
  INIT => X"0202000023022100"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10246_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12131\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2559\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1[7]_Z7235\: LUT6 
generic map(
  INIT => X"F0F1F0F1F1F1F3F3"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I1 => N_3811,
  I2 => N_3812,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.REEXCOVUV.UN18_LOCOV\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.REEXCOVUV.UN25_LOCOV\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.REEXCOVUV.UN13_LOCOV_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19[81]_Z7236\: LUT5 
generic map(
  INIT => X"CCF0AAF0"
)
port map (
  I0 => rfo1_data1(2),
  I1 => rfo2_data1(2),
  I2 => rfo2_data1(31),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(81));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19[76]_Z7237\: LUT5 
generic map(
  INIT => X"CFC0AFA0"
)
port map (
  I0 => rfo1_data1(7),
  I1 => rfo2_data1(7),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.OP1\(36),
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(76));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19[75]_Z7238\: LUT5 
generic map(
  INIT => X"FC0CFA0A"
)
port map (
  I0 => rfo1_data1(5),
  I1 => rfo2_data1(5),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.OP1\(40),
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(75));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19[73]_Z7239\: LUT6 
generic map(
  INIT => X"FF00F0F0CCCCAAAA"
)
port map (
  I0 => rfo1_data1(7),
  I1 => rfo1_data1(10),
  I2 => rfo2_data1(7),
  I3 => rfo2_data1(10),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I5 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(73));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19[72]_Z7240\: LUT5 
generic map(
  INIT => X"CFC0AFA0"
)
port map (
  I0 => rfo1_data1(11),
  I1 => rfo2_data1(11),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.OP1\(40),
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(72));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19[71]_Z7241\: LUT5 
generic map(
  INIT => X"FC0CFA0A"
)
port map (
  I0 => rfo1_data1(9),
  I1 => rfo2_data1(9),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.OP1\(44),
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(71));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19[69]_Z7242\: LUT6 
generic map(
  INIT => X"FF00F0F0CCCCAAAA"
)
port map (
  I0 => rfo1_data1(11),
  I1 => rfo1_data1(14),
  I2 => rfo2_data1(11),
  I3 => rfo2_data1(14),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I5 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(69));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19[66]_Z7243\: LUT5 
generic map(
  INIT => X"FC0CFA0A"
)
port map (
  I0 => rfo1_data1(14),
  I1 => rfo2_data1(14),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.OP1\(49),
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(66));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19[64]_Z7244\: LUT5 
generic map(
  INIT => X"FC0CFA0A"
)
port map (
  I0 => rfo1_data1(16),
  I1 => rfo2_data1(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.OP1\(51),
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(64));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41[254]_Z7245\: LUT6 
generic map(
  INIT => X"FF00F0F0CCCCAAAA"
)
port map (
  I0 => rfo1_data1(23),
  I1 => rfo1_data1(26),
  I2 => rfo2_data1(23),
  I3 => rfo2_data1(26),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I5 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41\(254));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41[253]_Z7246\: LUT6 
generic map(
  INIT => X"FF00F0F0CCCCAAAA"
)
port map (
  I0 => rfo1_data1(24),
  I1 => rfo1_data1(27),
  I2 => rfo2_data1(24),
  I3 => rfo2_data1(27),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I5 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41\(253));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[31]\: LUT6 
generic map(
  INIT => X"333355550F0F00FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8224\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[27]\: LUT6 
generic map(
  INIT => X"33330F0F00FF5555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8228\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A8[62]\: LUT6 
generic map(
  INIT => X"CC00CC0000000400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_722\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1344\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_776\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10948\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10925\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1[4]_Z7250\: LUT6 
generic map(
  INIT => X"FF7FFFFF00000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(254),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(253),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(256),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN4_NOTBINFNAN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTBINFNAN_0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1_0\(4),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1[3]_Z7251\: LUT5 
generic map(
  INIT => X"00151515"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(233),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN3_NOTAZERODENORM\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTAINFNAN_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTAINFNAN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[21]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF1F0F1100"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_741\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10246_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2764\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2214\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(21));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.EXTEND.TEMP[0]\: LUT6 
generic map(
  INIT => X"FFFEFFFAFFFEFFAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN26_XZYBUSLSBS\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN17_XZXBUS\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.EXTEND.TEMP[1]\: LUT5 
generic map(
  INIT => X"FFFFEAC0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.EXTEND.TEMP_0\(1),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN17_XZXBUS\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_I_A2[0]\: LUT6 
generic map(
  INIT => X"0080000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_I_A2_2\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_I_A2_1\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_I_A2_0\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_6\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_I_A2_3\(0),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_I_A2_4\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1101\);
\GRLFPC20.COMB.UN1_R.I.V_LUT6_2_RNIADOI1\: LUT6 
generic map(
  INIT => X"00FFCCFF00FFEFFF"
)
port map (
  I0 => \GRLFPC20.R.E.FPOP\,
  I1 => \GRLFPC20.R.M.FPOP\,
  I2 => \GRLFPC20.N_1538\,
  I3 => \GRLFPC20.N_1502_1\,
  I4 => \GRLFPC20.N_1536\,
  I5 => \GRLFPC20.N_1537\,
  O => \GRLFPC20.N_1494\);
\GRLFPC20.COMB.V.STATE14\: LUT6 
generic map(
  INIT => X"AAA8AAAA00000000"
)
port map (
  I0 => \GRLFPC20.R.I.V\,
  I1 => \GRLFPC20.N_1306\,
  I2 => \GRLFPC20.N_1307\,
  I3 => \GRLFPC20.N_1310\,
  I4 => \GRLFPC20.COMB.UN1_MEXC_1_0\,
  I5 => \GRLFPC20.COMB.V.I.EXEC_5\,
  O => \GRLFPC20.N_2000\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[40]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFF444F000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2229_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2601\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2602\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1192\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2230\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(40));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15[15]\: LUT6 
generic map(
  INIT => X"FFFFFFFFA0A0B3A0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_0\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_766\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2800\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2591\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_222\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2448\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1725\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_21_0_1_TZ[40]_Z7260\: LUT6 
generic map(
  INIT => X"FFFFFFFFAAAE000C"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1230\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1580\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_720\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12131\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1347\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2233\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_21_0_1_TZ\(40));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2[61]_Z7261\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF1700"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10693_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10893\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10882\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2\(61));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3[18]_Z7262\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF1000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_749\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2693\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9558_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1036\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9726\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3\(18));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_1[18]_Z7263\: LUT6_L 
generic map(
  INIT => X"222200002F220F00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9596\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_746\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9629\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9969_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_314_I\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12131\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_1\(18));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0[25]_Z7264\: LUT6 
generic map(
  INIT => X"FFFF000800080008"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12132\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9605_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9338_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12196_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9858_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_6_1\(25),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(25));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_0[25]_Z7265\: LUT6 
generic map(
  INIT => X"BAAAAAAA30000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_0_0\(25),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9366_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9605_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9338_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9389_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9709\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_0\(25));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2[34]_Z7266\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF0400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9366_I\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9739_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9967\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12180\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2\(34));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0[0]_Z7267\: LUT6_L 
generic map(
  INIT => X"3030220000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9723_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9338_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9666_1_I_0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0[35]_Z7268\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF0F1F0011"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9785_1_I_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_135\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12131\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_765\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1283\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0_0\(35),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(35));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15_1[16]_Z7269\: LUT6 
generic map(
  INIT => X"FFFFFFFF005000DC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1580\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2594\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_720\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12131\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2255\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15_1\(16));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_0[29]_Z7270\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFDC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_765\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2818\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1283\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2335\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2336\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2337\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_0\(29));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3[36]_Z7271\: LUT6 
generic map(
  INIT => X"FFFFFFFF0C004C00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_907\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9790_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10790\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10025_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_328\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0\(36),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3\(36));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0[36]_Z7272\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_76\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10006\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_328\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(36),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10023\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0\(36));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0[27]_Z7273\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF0009"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12132\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_398\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9779\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9799\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(27));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1[27]_Z7274\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_909\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9601_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10410\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9785\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9782\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(27));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2[13]_Z7275\: LUT4_L 
generic map(
  INIT => X"FFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10035\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9548\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9561\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9558\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2\(13));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3[13]_Z7276\: LUT6 
generic map(
  INIT => X"FEFAFCF0EEAACC00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_8_0\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_0_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_747_I\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_A2_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1234\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9551_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3\(13));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_1[13]_Z7277\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0100"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_776\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10332\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_741\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_775\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(13),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9549\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_1\(13));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4[53]_Z7278\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF1000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9946_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9389_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9604_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10290\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10297\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4\(53));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1[5]_Z7279\: LUT6 
generic map(
  INIT => X"FFFFFFFFF4F04400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_747_I\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12021_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2635\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_6095_A2_11_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2606\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_983\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[50]_Z7280\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF040404FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9887_I\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9671_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_717\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_742\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_765\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2150\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0\(50));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[44]_Z7281\: LUT6 
generic map(
  INIT => X"FFFFFFFFFF020202"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9700_I\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_369\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_921\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9324_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10030_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2210\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0\(44));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1[48]_Z7282\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF0800"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9576_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_261\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9738_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10158\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10156\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(48));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3[48]_Z7283\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9389_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9738_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9785_1_I_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10170\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10163\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3\(48));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1[55]_Z7284\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF0090"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9906_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_720\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10448\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10457\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(55));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2[55]_Z7285\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFD000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9657_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1149\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10765_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10449\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10442\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2\(55));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5[55]_Z7286\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0800"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10441_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1048_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9972_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9785_1_I_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_1\(55),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_966\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5\(55));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1[59]_Z7287\: LUT6_L 
generic map(
  INIT => X"CF0FCC00EFAFECA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A24_7_0\(59),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9642\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9969_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A24_0\(59),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A24_10_1\(59),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_775\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(59));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7[59]_Z7288\: LUT6 
generic map(
  INIT => X"FFFFFFFF08000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_52\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9604_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2600\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4\(59),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7\(59));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0[32]_Z7289\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF0080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9915_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9508_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9828\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_720\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9860\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(32),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(32));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0[32]_Z7290\: LUT6 
generic map(
  INIT => X"0040FFFF00400040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9840\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9338_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_1_1\(32),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0\(32));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_0[47]_Z7291\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0010"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_746\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12132\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9605_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_289\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10090\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_0_0\(47),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_0\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_5[47]_Z7292\: LUT6 
generic map(
  INIT => X"FFFFFFFFDFDD0F00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_314_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_715\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2605\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1002_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_5_0\(47),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_5\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_6_0[47]_Z7293\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_23_0\(47),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10790\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9394_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10088\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2_0\(47),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_3_0\(47),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_6_0\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_0[11]_Z7294\: LUT6 
generic map(
  INIT => X"FFFFFFFFFF040404"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9973_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_52\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9492_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_17_0\(11),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9326\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_0\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_6[11]_Z7295\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0032"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9505_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_125\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9558_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9785_1_I_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9316\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9318\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_6\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0[57]_Z7296\: LUT6 
generic map(
  INIT => X"FFFFFFFF80400000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9555_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10576\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9338_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(57),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1[57]_Z7297\: LUT6 
generic map(
  INIT => X"FFFFFFFFBAAA3000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_20_0\(57),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10592_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9605_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9972_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9558_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10616\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2[57]_Z7298\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF2020FF20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_6_0\(57),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9605_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1230\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10624_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10410\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10619\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6[57]_Z7299\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF0032"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10648\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10869\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10647\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_775\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9451\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_1\(57),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_1[57]_Z7300\: LUT6 
generic map(
  INIT => X"0000F1F000001100"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10640\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10654\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9969_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1019_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_304\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9670_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_1\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_6_1[31]_Z7301\: LUT6 
generic map(
  INIT => X"FFFFFFFF70007060"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9428\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9969_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10332\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_0\(31),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_6_1\(31));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_0[17]_Z7302\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0CAE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10895\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2591\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_742\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12131\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2447\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2448\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_0\(17));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7[19]_Z7303\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF8000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_759\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9338_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9972_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_967\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7_0\(19),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_1[19]_Z7304\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF02"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9915_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_304\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_720\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9660\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9661\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9663\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_1\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_1[33]_Z7305\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0010"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_59\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_304\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10410\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_720\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9928\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(33),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_1\(33));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7_0[33]_Z7306\: LUT6 
generic map(
  INIT => X"FFFFFFFFCC00ECA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9600_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9919_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1175\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1232\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_720\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0\(33),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7_0\(33));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3[52]_Z7307\: LUT6 
generic map(
  INIT => X"FFFFFFFF8080FF80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10236_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10888_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9861_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_9_1\(52),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0\(52),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6[54]_Z7308\: LUT6 
generic map(
  INIT => X"FFFFFFFFC0C0AA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_8_0\(54),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_741\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1272\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10948_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9394_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3\(54),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8_0[54]_Z7309\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF8000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9969_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9610_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10332\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1025\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0\(54),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8_0\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8_1[54]_Z7310\: LUT6 
generic map(
  INIT => X"BB00FBF0BB00BB00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_999_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10332\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1230\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_16_TZ\(54),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_775\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2724\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8_1\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9_0[54]_Z7311\: LUT5_L 
generic map(
  INIT => X"FFFFEAC0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2640\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10405\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10383_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2600\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_0\(54),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9_0\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_0[60]_Z7312\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF0800"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9946_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10790\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9652_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10090\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_0_1\(60),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_0\(60));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_4[60]_Z7313\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFE000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9577\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9790_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9601_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9972_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10824\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10839\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_4\(60));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_5[60]_Z7314\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0010"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12195\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9671_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_5_1\(60),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_534\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_5\(60));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2[56]_Z7315\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFF1F0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_906\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_796\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1012\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9670_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10535\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9604\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2\(56));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_6[56]_Z7316\: LUT6 
generic map(
  INIT => X"FFFFFFFF85000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9969_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_314_I\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9972_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_6_0\(56),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_6\(56));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIP48L1[91]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIR68L1[93]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIT88L1[93]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_3_Z7320\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(114),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN_1_Z7321\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIJ3BU[106]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIL5BU[107]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI0RJF[106]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIG0HF2[108]\: LUT5 
generic map(
  INIT => X"33A5FFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_812_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_515\);
\GRLFPC20.R.A.RF2REN_RNO_0[1]\: LUT3 
generic map(
  INIT => X"AC"
)
port map (
  I0 => cpi_d_inst(14),
  I1 => cpi_d_inst(25),
  I2 => \GRLFPC20.N_1583\,
  O => \GRLFPC20.N_2962\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI1TNQ1[86]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNICI0C1[86]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.UN84_TEMP_LUT6_2_RNINKV01\: LUT5 
generic map(
  INIT => X"CC5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.UN84_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIGM0C1[88]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.COMB.UN15_HOLDN_Z7331\: LUT4 
generic map(
  INIT => X"5A66"
)
port map (
  I0 => cpi_a_inst(7),
  I1 => rfo1_data2(31),
  I2 => rfo2_data2(31),
  I3 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.COMB.UN15_HOLDN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.UN348_TEMP_LUT6_2_RNIK32M1\: LUT5 
generic map(
  INIT => X"CC5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.UN348_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIJAJQ1[62]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3_Z7334\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_Z7335\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_2_Z7336\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_LUT6_2_RNIRG1V[6]\: LUT5 
generic map(
  INIT => X"CC5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.UN3_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIUVRB1[60]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_Z7339\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI02SB1[62]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI3F8L1[97]\: LUT5 
generic map(
  INIT => X"C3A5FFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_554\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI5H8L1[97]\: LUT5 
generic map(
  INIT => X"A5C3FFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_552\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI2VUB3[99]\: LUT5 
generic map(
  INIT => X"33A5FFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_803_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_550\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI75PO[100]\: LUT5 
generic map(
  INIT => X"A5C3FFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_544\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIB9PO[102]\: LUT5 
generic map(
  INIT => X"A5C3FFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_537\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIDBPO[103]\: LUT5 
generic map(
  INIT => X"A5C3FFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_523\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIFDPO[105]\: LUT5 
generic map(
  INIT => X"C3A5FFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_521\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIHFPO[105]\: LUT5 
generic map(
  INIT => X"A5C3FFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_519\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNINLPO[108]\: LUT5 
generic map(
  INIT => X"A5C3FFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_513\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIGFQO[110]\: LUT5 
generic map(
  INIT => X"C3A5FFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_499\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI99RO[110]\: LUT5 
generic map(
  INIT => X"A5C3FFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_457\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIBBRO[111]\: LUT5 
generic map(
  INIT => X"A5C3FFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_453\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1_Z7353\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(114),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_2_Z7354\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(114),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIOKLF[111]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIDDRO[113]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIMILF[110]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIDVCU[113]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNITOKF[110]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIBTCU[111]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIPRLQ[113]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI4VJF[108]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI9RCU[110]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNINPLQ[111]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI2TJF[107]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIG1CU[110]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNILNLQ[110]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI9PAU[101]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI7NAU[100]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI7EIC1[99]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIGO2C1[97]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.UN348_TEMP_LUT6_2_RNIVH5M1\: LUT5 
generic map(
  INIT => X"CC5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.UN462_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.UN18_TEMP_LUT6_2_RNIFDGB1\: LUT5 
generic map(
  INIT => X"CC5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.UN111_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNICK2C1[94]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI31QQ1[97]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIHV2N1[97]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIAI2C1[93]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIVA8L1[94]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI1VPQ1[95]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIFT2N1[97]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI8G2C1[93]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIVSPQ1[94]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIDR2N1[95]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI6E2C1[91]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIBP2N1[94]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI4C2C1[91]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIROPQ1[93]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI9N2N1[93]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIBI1C1[89]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIPMPQ1[91]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI7L2N1[93]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIIO0C1[88]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIU87L1[89]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNINKPQ1[91]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI3H2N1[91]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI3D6L1[88]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI51OQ1[88]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIAN1N1[89]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI3VNQ1[88]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIHT0N1[88]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIAG0C1[84]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIFR0N1[88]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI8E0C1[84]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIT66L1[84]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIVQNQ1[86]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIDP0N1[86]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI6C0C1[83]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIR46L1[84]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNITONQ1[84]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIBN0N1[86]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIP26L1[83]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIRMNQ1[84]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI9L0N1[84]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI17NT2[82]\: LUT5 
generic map(
  INIT => X"CC5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_846_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNILU5L1[80]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNININQ1[81]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI5H0N1[83]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNILGNQ1[80]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI3F0N1[81]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI3B4L1[78]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNISMMQ1[80]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI1D0N1[80]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI194L1[77]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI8JVM1[80]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIV64L1[76]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI1RLQ1[77]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIFPUM1[78]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIT44L1[75]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIVOLQ1[76]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIDNUM1[77]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI6AUB1[73]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_LUT6_2_RNIHTPD1[2]\: LUT5 
generic map(
  INIT => X"CC5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.UN393_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIBLUM1[76]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI48UB1[72]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIP04L1[73]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI26UB1[71]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIQKSB3[73]\: LUT5 
generic map(
  INIT => X"CC5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.UN213_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIPILQ1[73]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI7HUM1[75]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.UN36_TEMP_LUT6_2_RNIB5PT\: LUT5 
generic map(
  INIT => X"CC5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.UN36_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNILS3L1[71]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNINGLQ1[72]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI5FUM1[73]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI7ATB1[70]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIJQ3L1[70]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNILELQ1[71]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.UN555_TEMP_LUT6_2_RNI05MJ1\: LUT5 
generic map(
  INIT => X"CC5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.UN555_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIEGSB1[68]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIQ03L1[70]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIJCLQ1[70]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNICESB1[67]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIQIKQ1[70]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIACSB1[66]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI1PJQ1[68]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI8ASB1[66]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.UN18_TEMP_LUT6_2_RNIB6DB1\: LUT5 
generic map(
  INIT => X"CC5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.UN18_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNITKJQ1[66]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIBJSM1[67]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI46SB1[64]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.UN537_TEMP_LUT6_2_RNI9B3I1\: LUT5 
generic map(
  INIT => X"CC5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.UN537_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI24SB1[62]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIPGJQ1[64]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.UN537_TEMP_LUT6_2_RNIGNR21\: LUT4 
generic map(
  INIT => X"CA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.UN537_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.UN534_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_T_3[0]_Z7464\: LUT5 
generic map(
  INIT => X"AA91AA9D"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(377),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(375),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(376),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(374),
  I4 => N_3882,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_T_3\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_1_Z7465\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_2_Z7466\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIUOJF[105]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI34KQ[108]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.UN84_TEMP_LUT6_2_RNIU5PI\: LUT5 
generic map(
  INIT => X"CC5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.UN138_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI12KQ[107]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIH1BU[105]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIVVJQ[106]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIOIJF[102]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIFVAU[105]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNITTJQ[105]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIMGJF[101]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIDTAU[103]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIRRJQ[105]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIKEJF[100]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIBRAU[102]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIPPJQ[103]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIK5RT[99]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNINNJQ[102]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIKS2C1[99]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNILLJQ[101]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIIQ2C1[97]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.UN639_TEMP_LUT6_2_RNIAO481\: LUT5 
generic map(
  INIT => X"CC5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.UN639_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI4A0C1[81]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.UN36_TEMP_LUT6_2_RNIC7QT\: LUT5 
generic map(
  INIT => X"CC5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.UN66_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI9EVB1[80]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIGKUB1[78]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIEIUB1[77]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNICGUB1[76]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIAEUB1[75]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI8CUB1[75]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.UN198_TEMP_RNI51CF1\: LUT5 
generic map(
  INIT => X"CC5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.UN198_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIR02L1[66]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIPU1L1[64]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNINS1L1[64]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNILQ1L1[62]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNINEJQ1[64]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.UN180_TEMP_LUT6_2_RNIE9FJ1\: LUT5 
generic map(
  INIT => X"CC5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.UN180_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIHM1L1[60]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI19SM1[62]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIOS0L1[60]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_Z7506\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(114),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0[48]_Z7507\: LUT6_L 
generic map(
  INIT => X"00000303AA00AB03"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_7_0\(48),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_261\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9629\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9652_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_717\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(48));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR_0_Z7508\: LUT5 
generic map(
  INIT => X"000F1111"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR_1_Z7509\: LUT5 
generic map(
  INIT => X"00330505"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M12[1]_Z7510\: LUT5 
generic map(
  INIT => X"55445545"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_SS0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M12\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M12[0]_Z7511\: LUT6 
generic map(
  INIT => X"BBAABBABBBABBBAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_7\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_SS0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M12\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M12[2]_Z7512\: LUT6 
generic map(
  INIT => X"0000030200000303"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_SS0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M12\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15[17]\: LUT6 
generic map(
  INIT => X"AA000000AB030303"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9366_I\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9700_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_369\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9604_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2583\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_222\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1648\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15_2[17]\: LUT6 
generic map(
  INIT => X"F0000000F8888888"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1171\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9560_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9506_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9394_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12131\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1711\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_10[75]\: LUT6_L 
generic map(
  INIT => X"BEBB9C9936331411"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(51),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(52),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS\,
  I4 => N_3881,
  I5 => N_3882,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8814\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_14[142]_Z7516\: LUT6_L 
generic map(
  INIT => X"03AA00AAFCAA00AA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(144),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(376),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(374),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I5 => N_3882,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_14\(142));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9[57]_Z7517\: LUT6 
generic map(
  INIT => X"88000000A8A00000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10654\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9911_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1019_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1230\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10410\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9\(57));
\GRLFPC20.COMB.UN9_CCV_2_RNIOKQ21\: LUT5 
generic map(
  INIT => X"00151515"
)
port map (
  I0 => \GRLFPC20.COMB.UN9_CCV_2\,
  I1 => \GRLFPC20.R.I.EXEC\,
  I2 => \GRLFPC20.R.I.INST\(19),
  I3 => \GRLFPC20.R.X.AFSR\,
  I4 => \GRLFPC20.R.X.LD\,
  O => cpo_ccv);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A14_2[34]\: LUT6 
generic map(
  INIT => X"1104000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12021_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1230\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9967\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_A26[31]\: LUT6 
generic map(
  INIT => X"8A00880002000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9850_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1175\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9385\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13[25]\: LUT6 
generic map(
  INIT => X"0000000011150005"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_732\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12132\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9840\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_0\(11),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9716\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_1_A2[37]\: LUT6 
generic map(
  INIT => X"0000000000005004"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_746\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_741\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_969\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.TEMP_1_Z7523\: LUT6 
generic map(
  INIT => X"00000000AA22A022"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(73),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(74),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(71),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(75),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN10_S_MOV\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.TEMP_1\);
\GRLFPC20.RS1V_0_SQMUXA_0_A2\: LUT6 
generic map(
  INIT => X"0900000000000000"
)
port map (
  I0 => cpi_d_inst(19),
  I1 => cpi_d_inst(20),
  I2 => cpi_d_inst(23),
  I3 => cpi_d_inst(30),
  I4 => cpi_d_inst(31),
  I5 => \GRLFPC20.N_3109\,
  O => \GRLFPC20.RS1V_0_SQMUXA\);
\GRLFPC20.MOV_5_SQMUXA_0_A2_0\: LUT6 
generic map(
  INIT => X"0010000000000000"
)
port map (
  I0 => cpi_d_inst(19),
  I1 => cpi_d_inst(20),
  I2 => cpi_d_inst(23),
  I3 => cpi_d_inst(30),
  I4 => cpi_d_inst(31),
  I5 => \GRLFPC20.N_3109\,
  O => \GRLFPC20.N_3129\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN1_S_14_Z7526\: LUT5 
generic map(
  INIT => X"FFFCEEB7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN1_S_14\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_I_18_0_Z7527\: LUT6_L 
generic map(
  INIT => X"810F4200240018F0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(233),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(234),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1323\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(11),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(10),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_I_18_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0[30]_Z7528\: LUT5_L 
generic map(
  INIT => X"00F088F8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1333\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10891_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_222\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_765\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(30));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_1[26]_Z7529\: LUT6_L 
generic map(
  INIT => X"0F8F008800880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1170\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1561\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_751_I\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_328\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9669_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_1\(26));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0[36]_Z7530\: LUT6_L 
generic map(
  INIT => X"8888888F88888888"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_759\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_1_1\(36),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10948_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_328\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10410\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0\(36));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0[27]_Z7531\: LUT6 
generic map(
  INIT => X"FFFFFFFF00000054"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1229\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10006\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_909\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9786\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0\(27));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_0[53]_Z7532\: LUT6_L 
generic map(
  INIT => X"0F1F0F0F00110000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1048_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12132\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9506_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9558_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10948_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10690\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_0\(53));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0[4]_Z7533\: LUT6_L 
generic map(
  INIT => X"E0E0F9E000009900"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_0\(4),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10161_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_289\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10948_1\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_0[4]_Z7534\: LUT6_L 
generic map(
  INIT => X"88880000F888F000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10671_I\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9858_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9670_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10948_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10223_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_143\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_0\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1[28]_Z7535\: LUT6_L 
generic map(
  INIT => X"20200000FF20FF00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9461_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10584_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10948_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2823\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_765\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(28));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_0[5]_Z7536\: LUT6 
generic map(
  INIT => X"880088008800F8F0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_11378\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_2_0\(5),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10948_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2724\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_143\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_720\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_0\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0[7]_Z7537\: LUT6_L 
generic map(
  INIT => X"F0F00000F8F08800"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10869\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9558_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_157_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_1_1\(7),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_1[55]_Z7538\: LUT6 
generic map(
  INIT => X"ECDCCCCCA0500000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_9_0\(55),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9605_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10888_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10860\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10626_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_1\(55));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0[59]_Z7539\: LUT6 
generic map(
  INIT => X"CC00CC00CC00CDCD"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9549_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_831\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A24_19_1\(59),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9666_1_I_0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0\(59));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0[59]_Z7540\: LUT6 
generic map(
  INIT => X"4040FF400000FF00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10824_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_830\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_16_0\(52),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_715\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0\(59));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0[32]_Z7541\: LUT6_L 
generic map(
  INIT => X"F0F0F0F200000022"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9968_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9828\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9850_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9610_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_906\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_3_1\(32),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(32));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_0_0[47]_Z7542\: LUT6_L 
generic map(
  INIT => X"C0C00000D5C05500"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10734\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_766\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1344\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9667_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10087_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10790\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_0_0\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_6_1[47]_Z7543\: LUT6 
generic map(
  INIT => X"AAEAFFFF00C000C0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10767_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_9_0\(47),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2693\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9558_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9785_1_I_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2724\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_6_1\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2[11]_Z7544\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF73505050"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_59\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_831\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9330_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12021_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9652_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_13\(11),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_4_0[11]_Z7545\: LUT6 
generic map(
  INIT => X"F0001000F0000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_747_I\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9324_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_4_0\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0[57]_Z7546\: LUT6_L 
generic map(
  INIT => X"FF00FF4000004040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9505_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9605_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9969_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1230\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_9_1\(57),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_1[57]_Z7547\: LUT6 
generic map(
  INIT => X"AFAFAFAF00000020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9911_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_715\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9551_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_1\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_1[57]_Z7548\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFB9000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1229\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9666_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10891\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_1\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_5[31]_Z7549\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10332\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10888_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10025_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9394_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_991_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_5_1\(31),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_5\(31));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_2_0[31]_Z7550\: LUT6_L 
generic map(
  INIT => X"5F5F00005F5F0011"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_205\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1132_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_906\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10888_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_17_0\(11),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9666_1_I_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_2_0\(31));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_3_0[31]_Z7551\: LUT6_L 
generic map(
  INIT => X"D1111111C0000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_830\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9828\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_406\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9969_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9389_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_3_0\(31));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0[6]_Z7552\: LUT6_L 
generic map(
  INIT => X"F0F4F0FC004400CC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9490_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9748\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_143\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_720\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_0[19]_Z7553\: LUT6 
generic map(
  INIT => X"A0A0BBAAA0A0AAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_11_0\(19),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_783\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9604_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9738_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_717\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_0\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4[33]_Z7554\: LUT6_L 
generic map(
  INIT => X"DD5DCC0CCC0CCC0C"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_16\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9941\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12196_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9916_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10025_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1232\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4\(33));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_0[33]_Z7555\: LUT6 
generic map(
  INIT => X"30003A0A30003000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9739_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9508_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_234\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_A2_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10025_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_0\(33));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_0[24]_Z7556\: LUT6 
generic map(
  INIT => X"808080808080FF80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10948_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_157_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9861_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10943\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_765\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_0\(24));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0[52]_Z7557\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFFF01"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_411\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10584_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_795\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10225\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10767\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10237\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0[52]_Z7558\: LUT6_L 
generic map(
  INIT => X"88F8888800F00000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_6_0\(52),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1048_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A12_0\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_291_I\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9394_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9861_2\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_1[52]_Z7559\: LUT6_L 
generic map(
  INIT => X"C0EAC0C000AA0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_11_0\(52),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_7_0\(52),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9850_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10211\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9394_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9861_2\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_1\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_0[52]_Z7560\: LUT6 
generic map(
  INIT => X"FFFFFFFF0000AE0C"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9320_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9610_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_409\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9604_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_715\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10224\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_0\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0[54]_Z7561\: LUT6_L 
generic map(
  INIT => X"0000C0C00088C0C8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9637_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10405\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_234\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_795\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_289\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_0[54]_Z7562\: LUT6 
generic map(
  INIT => X"F0F0F8F000008800"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9600_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1019_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9389_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_906\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_22_0\(54),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_0\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_1[54]_Z7563\: LUT6 
generic map(
  INIT => X"808080808080FF80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9850_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1267\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_291_I\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9738_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9785_1_I_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_720\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_1\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_3[60]_Z7564\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF2010"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9739_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10819\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10827\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_3\(60));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_1_0[60]_Z7565\: LUT6 
generic map(
  INIT => X"FF000000FF101010"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_907\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9994_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9788_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A26_22_0\(60),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9785_1_I_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_1_0\(60));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_0[49]_Z7566\: LUT6 
generic map(
  INIT => X"BAAA300030003000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10592_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2162_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9972_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9671_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2606\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_0\(49));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_2[49]_Z7567\: LUT5 
generic map(
  INIT => X"FFFFFF10"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_254\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2591\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1041\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2166\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_2\(49));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_3[56]_Z7568\: LUT6 
generic map(
  INIT => X"FFFFFFFF33330020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10207_I_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1347\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10522\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_3\(56));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0[51]_Z7569\: LUT6_L 
generic map(
  INIT => X"22220000F222F000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_722\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_398\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9911_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1230\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9670_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12131\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(51));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_0[51]_Z7570\: LUT6_L 
generic map(
  INIT => X"01010000AB01AA00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_775\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_157_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2630\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_742\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_0\(51));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[10]\: LUT5 
generic map(
  INIT => X"555503F3"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_Z7572\: LUT6 
generic map(
  INIT => X"53F35FFFFFAFFCAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[4]\: LUT5 
generic map(
  INIT => X"3333505F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(238),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(53));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS[9]_Z7574\: LUT6 
generic map(
  INIT => X"20202020E0202020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(235),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(9));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS[8]_Z7575\: LUT6 
generic map(
  INIT => X"20202020E0202020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(236),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(8));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[2]\: LUT5 
generic map(
  INIT => X"3333505F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(12),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(55));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[6]\: LUT5 
generic map(
  INIT => X"3333505F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(240),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(51));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[25]\: LUT6 
generic map(
  INIT => X"333327270F332727"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(32));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[5]\: LUT5 
generic map(
  INIT => X"3333505F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(239),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[7]\: LUT5 
generic map(
  INIT => X"3333505F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(241),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(50));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[12]\: LUT6 
generic map(
  INIT => X"5555535333555353"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(45));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[33]\: LUT6 
generic map(
  INIT => X"0F0F1D1D550F1D1D"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(24));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[22]\: LUT6 
generic map(
  INIT => X"5555535333555353"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(35));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[26]\: LUT6 
generic map(
  INIT => X"3333353555333535"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(31));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[13]\: LUT6 
generic map(
  INIT => X"5555535333555353"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(44));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[37]\: LUT6 
generic map(
  INIT => X"5555535333555353"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(20));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[15]\: LUT6 
generic map(
  INIT => X"5555535333555353"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(42));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[11]\: LUT6 
generic map(
  INIT => X"5555535333555353"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(46));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[8]\: LUT5 
generic map(
  INIT => X"3333505F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(242),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(49));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[14]\: LUT6 
generic map(
  INIT => X"5555535333555353"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(43));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[30]\: LUT6 
generic map(
  INIT => X"3333353555333535"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(27));
\GRLFPC20.FPI.OP2[34]_Z7592\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(2),
  I1 => rfo2_data2(2),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(34));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_Z7593\: LUT6 
generic map(
  INIT => X"5F5F33FFFAFAFFCC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[38]\: LUT6 
generic map(
  INIT => X"5555535333555353"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[35]\: LUT6 
generic map(
  INIT => X"5555535333555353"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(22));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[34]\: LUT6 
generic map(
  INIT => X"5555535333555353"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(23));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[16]\: LUT6 
generic map(
  INIT => X"5555535333555353"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(41));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[377]\: LUT5_L 
generic map(
  INIT => X"0010FFBF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(5),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I4 => N_3880,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_I\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[31]\: LUT6 
generic map(
  INIT => X"0F0F1D1D550F1D1D"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(26));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[29]\: LUT6 
generic map(
  INIT => X"0F0F1D1D550F1D1D"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(28));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0[3]\: LUT5 
generic map(
  INIT => X"3333505F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(237),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_0_CY_RNO\: LUT6 
generic map(
  INIT => X"8F88FFF807007770"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(5),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8372\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN8_TEMP\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_I_29\: LUT6 
generic map(
  INIT => X"E0201FDF1FDFE020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(240),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(4),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12032\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A15_2[18]\: LUT6 
generic map(
  INIT => X"00000000880A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9601_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_796\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9601\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A14_4[34]\: LUT6 
generic map(
  INIT => X"D080000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9969_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9969_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9969\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_4[55]\: LUT6_L 
generic map(
  INIT => X"0000000013020000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1230\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_775\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10442\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_1[61]\: LUT6_L 
generic map(
  INIT => X"00000000B0100000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9461_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_304\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10884\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2_1[60]_Z7608\: LUT6 
generic map(
  INIT => X"FFFFFFFF00008D00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9404_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_715\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10834\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2_1\(60));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS_1_0[7]\: LUT6 
generic map(
  INIT => X"20202020E0202020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(237),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M13[0]_Z7610\: LUT5 
generic map(
  INIT => X"BABAFF00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_7_REP1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_8_REP1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_9_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_SS9\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_9\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M13\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1_Z7611\: LUT5 
generic map(
  INIT => X"88888880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(10),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(11),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN12_SRTOSTICKY_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_14[172]_Z7612\: LUT5_L 
generic map(
  INIT => X"01000E00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(376),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(374),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => N_3882,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_14\(172));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_12_Z7613\: LUT6 
generic map(
  INIT => X"965AF05A3CF05AF0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(232),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(245),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1323\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_12\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_I_36\: LUT6 
generic map(
  INIT => X"965AF05A3CF05AF0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(232),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(245),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1323\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12030\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1[5]_Z7615\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(241),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(243),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(240),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1_0\(5),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN3_NOTAZERODENORM\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_0[48]\: LUT6_L 
generic map(
  INIT => X"590A000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9508_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9738_1\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10155\);
\GRLFPC20.COMB.UN2_HOLDN\: LUT5 
generic map(
  INIT => X"10000000"
)
port map (
  I0 => cpi_a_annul,
  I1 => cpi_a_trap,
  I2 => holdn,
  I3 => \GRLFPC20.R.A.MOV\,
  I4 => \GRLFPC20.R.A.FPOP\,
  O => \GRLFPC20.N_1858\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN10_S_MOV_Z7618\: LUT6 
generic map(
  INIT => X"0100000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9490_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_234\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN10_S_MOV\);
\GRLFPC20.COMB.UN19_IUEXEC\: LUT5 
generic map(
  INIT => X"00020000"
)
port map (
  I0 => \GRLFPC20.R.MK.BUSY2\,
  I1 => \GRLFPC20.R.MK.BUSY\,
  I2 => \GRLFPC20.R.MK.RST\,
  I3 => \GRLFPC20.R.MK.RST2\,
  I4 => \GRLFPC20.N_2103\,
  O => \GRLFPC20.N_2102\);
\GRLFPC20.COMB.SEQERR.UN3_QNE_1\: LUT5 
generic map(
  INIT => X"00040000"
)
port map (
  I0 => cpi_d_inst(19),
  I1 => cpi_d_inst(20),
  I2 => cpi_d_inst(22),
  I3 => cpi_d_inst(23),
  I4 => \GRLFPC20.COMB.SEQERR.UN3_QNE_1_0\,
  O => \GRLFPC20.COMB.V.A.AFQ_1_1\);
\GRLFPC20.RS2_0_SQMUXA\: LUT6 
generic map(
  INIT => X"0400000000000000"
)
port map (
  I0 => cpi_d_inst(20),
  I1 => cpi_d_inst(21),
  I2 => cpi_d_inst(22),
  I3 => cpi_d_inst(23),
  I4 => cpi_d_inst(24),
  I5 => \GRLFPC20.N_878\,
  O => \GRLFPC20.N_1583\);
\GRLFPC20.COMB.RDD_1.M4_E_I_A3_0\: LUT6 
generic map(
  INIT => X"0010000000000000"
)
port map (
  I0 => cpi_d_inst(6),
  I1 => cpi_d_inst(9),
  I2 => cpi_d_inst(12),
  I3 => cpi_d_inst(13),
  I4 => \GRLFPC20.N_3117\,
  I5 => \GRLFPC20.N_3123\,
  O => \GRLFPC20.N_3084\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A8_3[62]\: LUT6 
generic map(
  INIT => X"0000000A0000002A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_76\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_831\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_776\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12195\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10929\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3[54]_Z7624\: LUT6_L 
generic map(
  INIT => X"0000000080008202"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9490_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_795\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_328\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTAINFNAN_2_Z7625\: LUT6_L 
generic map(
  INIT => X"C0008000C0000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(234),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(241),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(240),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN8_NOTAINFNAN_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTAINFNAN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.EXTEND.TEMP_0[1]_Z7626\: LUT5_L 
generic map(
  INIT => X"EAAAC000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(230),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(11),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.EXTEND.TEMP_0\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_0[61]_Z7627\: LUT6 
generic map(
  INIT => X"FF80008000800080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9461_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_76\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9969_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9911_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_5_0\(48),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9558_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_0\(61));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0[18]_Z7628\: LUT6_L 
generic map(
  INIT => X"00002222A000A222"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9994_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9629\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_749\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9969_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10332\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_741\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0\(18));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0[34]_Z7629\: LUT6_L 
generic map(
  INIT => X"30003000BAAA3000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9975_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10332\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9652_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10025_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9738_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(34));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0_0[35]_Z7630\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF00009000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_291_I\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9394_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_720\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2233\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0_0\(35));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0[36]_Z7631\: LUT6 
generic map(
  INIT => X"0000808000CC80CC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_768_I\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_205\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_783\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10410\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(36));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_0[5]_Z7632\: LUT6 
generic map(
  INIT => X"04040404FF040404"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1331\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_749\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9671_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1333\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9861_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_0\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0[59]_Z7633\: LUT6_L 
generic map(
  INIT => X"3030703400004004"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10824_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_409\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10759_2\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0\(59));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_3_0[47]_Z7634\: LUT6_L 
generic map(
  INIT => X"F2F0220022002200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10767_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9667_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9605_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9911_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9601_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9652_1\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_3_0\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0[57]_Z7635\: LUT6_L 
generic map(
  INIT => X"CC40CC0040400000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10207_I_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1149\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10629_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10631_2\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_5_1[31]_Z7636\: LUT6_L 
generic map(
  INIT => X"1504000011000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1553_I\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9671_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10025_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9738_1\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_5_1\(31));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7_0[19]_Z7637\: LUT6_L 
generic map(
  INIT => X"00F000F000008888"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1132_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9664_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9972_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_717\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7_0\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0[33]_Z7638\: LUT6_L 
generic map(
  INIT => X"55D5008000800080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9600_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12021_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_796\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10888_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_17_0\(11),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0\(33));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0[54]_Z7639\: LUT6_L 
generic map(
  INIT => X"55550000D555C000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_211\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_768_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9850_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1019_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9738_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9666_1_I_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7_1[54]_Z7640\: LUT6_L 
generic map(
  INIT => X"C0EAC0C000AA0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_289\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10891_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_717\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10626_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7_1\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_1_0[56]_Z7641\: LUT6_L 
generic map(
  INIT => X"002200220022F0F2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9503_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_732\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_328\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9666_1_I_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10410\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_1_0\(56));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN11_WQSTSETS_0_Z7642\: LUT6 
generic map(
  INIT => X"F777F777F7770777"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(14),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(4),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(5),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN11_WQSTSETS_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0_0_0[0]_Z7643\: LUT6 
generic map(
  INIT => X"DFFF0000DF000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_30_REP1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_29_REP1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_FAST\(10),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0_0_0\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.RESULT_IV_0[1]_Z7644\: LUT6 
generic map(
  INIT => X"2AEAAAAA2A2AAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(59),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(49),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(51),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(52),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(50),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SFTLFT.AREGXORBREG\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.RESULT_IV_0\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_RNO[16]\: LUT4_L 
generic map(
  INIT => X"D515"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(16),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(4),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_870_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_RNO[14]\: LUT4_L 
generic map(
  INIT => X"15D5"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(16),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(5),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_871_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[33]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(21),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(149),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7884\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5[24]_Z7648\: LUT6 
generic map(
  INIT => X"33300300AAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(291),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(24));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[41]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(13),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(157),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7876\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[46]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(8),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(162),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7871\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[51]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(3),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(167),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7866\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5[57]_Z7652\: LUT6 
generic map(
  INIT => X"0F0C0300AAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(258),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS[6]_Z7653\: LUT5 
generic map(
  INIT => X"E0202020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(238),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS[5]_Z7654\: LUT5 
generic map(
  INIT => X"E0202020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(239),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M8[1]_Z7655\: LUT3_L 
generic map(
  INIT => X"54"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST\(7),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST\(9),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M8\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M13[2]_Z7656\: LUT5 
generic map(
  INIT => X"00110010"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_3_REP1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M8\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M13\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5[9]_Z7657\: LUT6 
generic map(
  INIT => X"33300300AAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(306),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(9));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[29]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(25),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(145),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7888\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5[55]_Z7659\: LUT6 
generic map(
  INIT => X"33003030AAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(260),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(55));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5[22]_Z7660\: LUT6 
generic map(
  INIT => X"33300300AAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(293),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(22));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5[21]_Z7661\: LUT6 
generic map(
  INIT => X"33003030AAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(294),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(21));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_6[75]\: LUT5 
generic map(
  INIT => X"AA695569"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(48),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(13),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(12),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(52),
  I4 => N_3812,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8810\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_1[5]\: LUT6 
generic map(
  INIT => X"33300300AAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(310),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[49]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(5),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(165),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7868\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[45]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(9),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(161),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7872\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_2[0]_Z7666\: LUT5 
generic map(
  INIT => X"CCCCD8CC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(5),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_2\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0[3]\: LUT5 
generic map(
  INIT => X"FFEF0040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(5),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I4 => \GRLFPC20.FPO.FRAC\(52),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0[2]\: LUT5 
generic map(
  INIT => X"FFEF0040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(5),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I4 => \GRLFPC20.FPO.FRAC\(53),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0[1]\: LUT5 
generic map(
  INIT => X"FFEF0040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(5),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I4 => \GRLFPC20.FPO.FRAC\(54),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0[0]\: LUT5 
generic map(
  INIT => X"FFEF0040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(5),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I4 => N_3880,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[52]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(2),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(168),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7865\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[50]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(4),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(166),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7867\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[48]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(6),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(164),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7869\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[47]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(7),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(163),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7870\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[44]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(10),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(160),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7873\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[43]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(11),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(159),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7874\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[42]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(12),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(158),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7875\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[39]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(155),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7878\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[38]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(16),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(154),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7879\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[37]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(17),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(153),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7880\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[36]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(18),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(152),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7881\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[35]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(19),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(151),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7882\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[34]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(20),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(150),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7883\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[32]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(22),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(148),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7885\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[30]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(24),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(146),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7887\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[28]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(26),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(144),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7889\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[27]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(27),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(143),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7890\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2[115]\: LUT5 
generic map(
  INIT => X"33B30080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(118),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => N_3825,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9071\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2[114]\: LUT5 
generic map(
  INIT => X"33B30080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(117),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
  I4 => N_3826,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9072\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5[7]_Z7690\: LUT6 
generic map(
  INIT => X"33300300AAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(308),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5[10]_Z7691\: LUT6 
generic map(
  INIT => X"33003030AAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(305),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(10));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5[14]_Z7692\: LUT6 
generic map(
  INIT => X"33300300AAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(301),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(14));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5[16]_Z7693\: LUT6 
generic map(
  INIT => X"33003030AAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(299),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(16));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5[18]_Z7694\: LUT6 
generic map(
  INIT => X"33003030AAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(297),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(18));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5[20]_Z7695\: LUT6 
generic map(
  INIT => X"33003030AAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(295),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(20));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5[27]_Z7696\: LUT6 
generic map(
  INIT => X"33003030AAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(288),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(27));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5[31]_Z7697\: LUT6 
generic map(
  INIT => X"33003030AAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(284),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(31));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5[40]_Z7698\: LUT6 
generic map(
  INIT => X"33003030AAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(275),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(40));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5[42]_Z7699\: LUT6 
generic map(
  INIT => X"33003030AAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(273),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(42));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5[45]_Z7700\: LUT6 
generic map(
  INIT => X"33300300AAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(270),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(45));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5[49]_Z7701\: LUT6 
generic map(
  INIT => X"33003030AAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(266),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(49));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M_RNO_1[2]\: LUT5_L 
generic map(
  INIT => X"2222222E"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(58),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\,
  I2 => \GRLFPC20.FPO.FRAC\(54),
  I3 => N_3881,
  I4 => N_3880,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.RESULT\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[54]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(170),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7863\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[53]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(169),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7864\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[40]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(14),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(156),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7877\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[31]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(23),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(147),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7886\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3[26]\: LUT4 
generic map(
  INIT => X"0ACC"
)
port map (
  I0 => rfo2_data2(28),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(142),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7891\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5[13]_Z7708\: LUT6 
generic map(
  INIT => X"33003030AAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(302),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(13));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5[35]_Z7709\: LUT6 
generic map(
  INIT => X"33003030AAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(280),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(35));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5[47]_Z7710\: LUT6 
generic map(
  INIT => X"33003030AAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(268),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5[2]_Z7711\: LUT6 
generic map(
  INIT => X"33300300AAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(313),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI073D1[41]\: LUT4_L 
generic map(
  INIT => X"A080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(41),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(38),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(39),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(40),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_591_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.EXPYBUS_1_I_A2_I[1]\: LUT3 
generic map(
  INIT => X"EA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(29),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(30),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_FAST\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_584\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3[1]_Z7714\: LUT5 
generic map(
  INIT => X"F0CCAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(372),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(1));
\GRLFPC20.COMB.DBGDATA_4[23]\: LUT5 
generic map(
  INIT => X"F3E2D1C0"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => \GRLFPC20.R.FSR.TEM\(0),
  I3 => rfo1_data1(23),
  I4 => rfo2_data1(23),
  O => cpo_dbg_data(23));
\GRLFPC20.COMB.UN1_FPCI_4_Z7716\: LUT5 
generic map(
  INIT => X"BA303030"
)
port map (
  I0 => cpi_a_cnt(1),
  I1 => \GRLFPC20.R.A.RS2D\,
  I2 => \GRLFPC20.R.A.RS2\(0),
  I3 => \GRLFPC20.R.A.RS1D\,
  I4 => \GRLFPC20.R.A.ST\,
  O => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20.COMB.UN1_R.A.RS1_1_Z7717\: LUT4 
generic map(
  INIT => X"AC0C"
)
port map (
  I0 => cpi_a_cnt(1),
  I1 => \GRLFPC20.R.A.RS1\(0),
  I2 => \GRLFPC20.R.A.RS1D\,
  I3 => \GRLFPC20.R.A.ST\,
  O => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20.COMB.DBGDATA_4[13]\: LUT6 
generic map(
  INIT => X"3F332E221D110C00"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => \GRLFPC20.R.STATE\(0),
  I3 => \GRLFPC20.R.STATE\(1),
  I4 => rfo1_data1(13),
  I5 => rfo2_data1(13),
  O => cpo_dbg_data(13));
\GRLFPC20.COMB.DBGDATA_4[25]\: LUT5 
generic map(
  INIT => X"F3E2D1C0"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => \GRLFPC20.R.FSR.TEM\(2),
  I3 => rfo1_data1(25),
  I4 => rfo2_data1(25),
  O => cpo_dbg_data(25));
\GRLFPC20.COMB.DBGDATA_4[16]\: LUT5 
generic map(
  INIT => X"F3E2D1C0"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => \GRLFPC20.R.FSR.FTT\(2),
  I3 => rfo1_data1(16),
  I4 => rfo2_data1(16),
  O => cpo_dbg_data(16));
\GRLFPC20.COMB.DBGDATA_4[24]\: LUT5 
generic map(
  INIT => X"F3E2D1C0"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => \GRLFPC20.R.FSR.TEM\(1),
  I3 => rfo1_data1(24),
  I4 => rfo2_data1(24),
  O => cpo_dbg_data(24));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1_I_0[3]\: LUT4 
generic map(
  INIT => X"05C5"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\);
\GRLFPC20.COMB.DBGDATA_4[31]\: LUT5 
generic map(
  INIT => X"F3E2D1C0"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => \GRLFPC20.R.FSR.RD\(1),
  I3 => rfo1_data1(31),
  I4 => rfo2_data1(31),
  O => cpo_dbg_data(31));
\GRLFPC20.COMB.DBGDATA_4[30]\: LUT5 
generic map(
  INIT => X"F3E2D1C0"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => \GRLFPC20.R.FSR.RD\(0),
  I3 => rfo1_data1(30),
  I4 => rfo2_data1(30),
  O => cpo_dbg_data(30));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2[247]\: LUT5_L 
generic map(
  INIT => X"BF8FB080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(234),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
  I3 => N_3811,
  I4 => \GRLFPC20.FPO.EXP\(10),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8788\);
\GRLFPC20.COMB.DBGDATA_4[10]\: LUT5 
generic map(
  INIT => X"F3E2D1C0"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => NN_1,
  I3 => rfo1_data1(10),
  I4 => rfo2_data1(10),
  O => cpo_dbg_data(10));
\GRLFPC20.COMB.DBGDATA_4[11]\: LUT5 
generic map(
  INIT => X"F3E2D1C0"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => CPO_CC_3,
  I3 => rfo1_data1(11),
  I4 => rfo2_data1(11),
  O => cpo_dbg_data(11));
\GRLFPC20.COMB.DBGDATA_4[14]\: LUT5 
generic map(
  INIT => X"F3E2D1C0"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => \GRLFPC20.R.FSR.FTT\(0),
  I3 => rfo1_data1(14),
  I4 => rfo2_data1(14),
  O => cpo_dbg_data(14));
\GRLFPC20.COMB.DBGDATA_4[0]\: LUT5 
generic map(
  INIT => X"F3E2D1C0"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => \GRLFPC20.R.FSR.CEXC\(0),
  I3 => rfo1_data1(0),
  I4 => rfo2_data1(0),
  O => cpo_dbg_data(0));
\GRLFPC20.COMB.DBGDATA_4[1]\: LUT5 
generic map(
  INIT => X"F3E2D1C0"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => \GRLFPC20.R.FSR.CEXC\(1),
  I3 => rfo1_data1(1),
  I4 => rfo2_data1(1),
  O => cpo_dbg_data(1));
\GRLFPC20.COMB.DBGDATA_4[2]\: LUT5 
generic map(
  INIT => X"F3E2D1C0"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => \GRLFPC20.R.FSR.CEXC\(2),
  I3 => rfo1_data1(2),
  I4 => rfo2_data1(2),
  O => cpo_dbg_data(2));
\GRLFPC20.COMB.DBGDATA_4[3]\: LUT5 
generic map(
  INIT => X"F3E2D1C0"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => \GRLFPC20.R.FSR.CEXC\(3),
  I3 => rfo1_data1(3),
  I4 => rfo2_data1(3),
  O => cpo_dbg_data(3));
\GRLFPC20.COMB.DBGDATA_4[4]\: LUT5 
generic map(
  INIT => X"F3E2D1C0"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => \GRLFPC20.R.FSR.CEXC\(4),
  I3 => rfo1_data1(4),
  I4 => rfo2_data1(4),
  O => cpo_dbg_data(4));
\GRLFPC20.COMB.DBGDATA_4[5]\: LUT5 
generic map(
  INIT => X"F3E2D1C0"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => \GRLFPC20.R.FSR.AEXC\(0),
  I3 => rfo1_data1(5),
  I4 => rfo2_data1(5),
  O => cpo_dbg_data(5));
\GRLFPC20.COMB.DBGDATA_4[6]\: LUT5 
generic map(
  INIT => X"F3E2D1C0"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => \GRLFPC20.R.FSR.AEXC\(1),
  I3 => rfo1_data1(6),
  I4 => rfo2_data1(6),
  O => cpo_dbg_data(6));
\GRLFPC20.COMB.DBGDATA_4[7]\: LUT5 
generic map(
  INIT => X"F3E2D1C0"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => \GRLFPC20.R.FSR.AEXC\(2),
  I3 => rfo1_data1(7),
  I4 => rfo2_data1(7),
  O => cpo_dbg_data(7));
\GRLFPC20.COMB.DBGDATA_4[8]\: LUT5 
generic map(
  INIT => X"F3E2D1C0"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => \GRLFPC20.R.FSR.AEXC\(3),
  I3 => rfo1_data1(8),
  I4 => rfo2_data1(8),
  O => cpo_dbg_data(8));
\GRLFPC20.COMB.DBGDATA_4[9]\: LUT5 
generic map(
  INIT => X"F3E2D1C0"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => \GRLFPC20.R.FSR.AEXC\(4),
  I3 => rfo1_data1(9),
  I4 => rfo2_data1(9),
  O => cpo_dbg_data(9));
\GRLFPC20.COMB.DBGDATA_4[15]\: LUT5 
generic map(
  INIT => X"F3E2D1C0"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => \GRLFPC20.R.FSR.FTT\(1),
  I3 => rfo1_data1(15),
  I4 => rfo2_data1(15),
  O => cpo_dbg_data(15));
\GRLFPC20.COMB.DBGDATA_4[22]\: LUT5 
generic map(
  INIT => X"F3E2D1C0"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => \GRLFPC20.R.FSR.NONSTD\,
  I3 => rfo1_data1(22),
  I4 => rfo2_data1(22),
  O => cpo_dbg_data(22));
\GRLFPC20.COMB.DBGDATA_4[26]\: LUT5 
generic map(
  INIT => X"F3E2D1C0"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => \GRLFPC20.R.FSR.TEM\(3),
  I3 => rfo1_data1(26),
  I4 => rfo2_data1(26),
  O => cpo_dbg_data(26));
\GRLFPC20.COMB.DBGDATA_4[27]\: LUT5 
generic map(
  INIT => X"F3E2D1C0"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => \GRLFPC20.R.FSR.TEM\(4),
  I3 => rfo1_data1(27),
  I4 => rfo2_data1(27),
  O => cpo_dbg_data(27));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1_I_0[0]\: LUT4 
generic map(
  INIT => X"90FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(257),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN26_XZYBUSLSBS_Z7744\: LUT5 
generic map(
  INIT => X"A888A000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(231),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(9),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(12),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(11),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(374),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN26_XZYBUSLSBS\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN8_TEMP_2[0]\: LUT6_L 
generic map(
  INIT => X"F7E6B3A2D5C49180"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_FAST\(10),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8372\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2[254]\: LUT5_L 
generic map(
  INIT => X"BFB08F80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(241),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
  I3 => \GRLFPC20.FPO.EXP\(3),
  I4 => \GRLFPC20.FPO.EXP\(4),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8781\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2[253]\: LUT5_L 
generic map(
  INIT => X"BFB08F80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(240),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
  I3 => \GRLFPC20.FPO.EXP\(4),
  I4 => \GRLFPC20.FPO.EXP\(5),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8782\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2[249]\: LUT5_L 
generic map(
  INIT => X"BFB08F80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(236),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
  I3 => \GRLFPC20.FPO.EXP\(8),
  I4 => \GRLFPC20.FPO.EXP\(9),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8786\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2[248]\: LUT5_L 
generic map(
  INIT => X"BFB08F80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(235),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
  I3 => \GRLFPC20.FPO.EXP\(9),
  I4 => \GRLFPC20.FPO.EXP\(10),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8787\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_Z7750\: LUT6 
generic map(
  INIT => X"EFEEAFAACFCC0F00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(13),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(375),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(16),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(9),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(11),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15[45]\: LUT6 
generic map(
  INIT => X"0000120000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(45));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_I_A2_0[0]_Z7752\: LUT6 
generic map(
  INIT => X"0000000000000013"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1186\);
\GRLFPC20.COMB.LOCKGEN.DEPCHECK\: LUT5 
generic map(
  INIT => X"FFFFFFFE"
)
port map (
  I0 => \GRLFPC20.R.A.FPOP\,
  I1 => \GRLFPC20.R.E.FPOP\,
  I2 => \GRLFPC20.R.M.FPOP\,
  I3 => \GRLFPC20.R.I.EXEC\,
  I4 => \GRLFPC20.R.X.FPOP\,
  O => \GRLFPC20.N_2103\);
\GRLFPC20.V.FSR.FTT_1_SQMUXA\: LUT6 
generic map(
  INIT => X"00000000F7F700F7"
)
port map (
  I0 => \GRLFPC20.R.X.AFQ\,
  I1 => \GRLFPC20.R.STATE\(1),
  I2 => \GRLFPC20.R.STATE\(0),
  I3 => \GRLFPC20.R.X.AFSR\,
  I4 => \GRLFPC20.R.X.LD\,
  I5 => \GRLFPC20.R.X.SEQERR\,
  O => \GRLFPC20.N_1421\);
\GRLFPC20.COMB.FPDECODE.ST_0_A2\: LUT6 
generic map(
  INIT => X"0200000000000000"
)
port map (
  I0 => cpi_d_inst(21),
  I1 => cpi_d_inst(22),
  I2 => cpi_d_inst(23),
  I3 => cpi_d_inst(24),
  I4 => cpi_d_inst(30),
  I5 => cpi_d_inst(31),
  O => \GRLFPC20.COMB.FPDECODE.ST\);
\GRLFPC20.COMB.FPDECODE.FPOP3\: LUT6 
generic map(
  INIT => X"0020000000000000"
)
port map (
  I0 => cpi_d_inst(19),
  I1 => cpi_d_inst(20),
  I2 => cpi_d_inst(21),
  I3 => cpi_d_inst(22),
  I4 => cpi_d_inst(23),
  I5 => cpi_d_inst(24),
  O => \GRLFPC20.N_940\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M14S2\: LUT5 
generic map(
  INIT => X"FFFEFFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_7_REP1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_8_REP1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_9_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_9\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_SM12\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD\: LUT6 
generic map(
  INIT => X"FEEEFCCCFAAAF000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST\(376),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(14),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(16),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(9),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(11),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\);
\GRLFPC20.COMB.UN9_CCV_2_Z7759\: LUT6 
generic map(
  INIT => X"FEFCFAF0EECCAA00"
)
port map (
  I0 => cpi_e_inst(19),
  I1 => cpi_m_inst(19),
  I2 => cpi_x_inst(19),
  I3 => \GRLFPC20.R.E.FPOP\,
  I4 => \GRLFPC20.R.M.FPOP\,
  I5 => \GRLFPC20.R.X.FPOP\,
  O => \GRLFPC20.COMB.UN9_CCV_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1_3[6]_Z7760\: LUT5 
generic map(
  INIT => X"FFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(250),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(251),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(252),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(257),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1_2\(6),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1_3\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTBINFNAN_0_Z7761\: LUT5 
generic map(
  INIT => X"80000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(250),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(251),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(252),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(255),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(257),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTBINFNAN_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_I_A2_0_2[0]\: LUT6 
generic map(
  INIT => X"0000000000000001"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_I_A2_0\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_I_A2_1_0[0]\: LUT6 
generic map(
  INIT => X"0000000000000001"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_I_A2_1\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_I_A2_2[0]_Z7764\: LUT6 
generic map(
  INIT => X"0000000000000001"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_I_A2_2\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_I_A2_3[0]_Z7765\: LUT6 
generic map(
  INIT => X"0000000000000001"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_I_A2_3\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN3_S_SQRT_0_Z7766\: LUT5 
generic map(
  INIT => X"00000100"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN3_S_SQRT_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_7_RNIQE402\: LUT6 
generic map(
  INIT => X"FFFFFFFEFFFFFFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST\(17),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_7\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_I_I_A2_0_O2_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0_0_O2_0[2]_Z7768\: LUT5 
generic map(
  INIT => X"EEF00000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_30_REP1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_29_REP1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(242),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0_0_O2_0\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_3_Z7769\: LUT5 
generic map(
  INIT => X"80000000"
)
port map (
  I0 => \GRLFPC20.FPO.FRAC\(47),
  I1 => \GRLFPC20.FPO.FRAC\(48),
  I2 => \GRLFPC20.FPO.FRAC\(49),
  I3 => \GRLFPC20.FPO.FRAC\(52),
  I4 => \GRLFPC20.FPO.FRAC\(53),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.REEXCOVUV.UN13_LOCOV_2_Z7770\: LUT6_L 
generic map(
  INIT => X"8000000000000000"
)
port map (
  I0 => \GRLFPC20.FPO.EXP\(1),
  I1 => \GRLFPC20.FPO.EXP\(2),
  I2 => \GRLFPC20.FPO.EXP\(3),
  I3 => \GRLFPC20.FPO.EXP\(4),
  I4 => \GRLFPC20.FPO.EXP\(7),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.REEXCOVUV.UN13_LOCOV_0_2\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.REEXCOVUV.UN13_LOCOV_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN30_CONDITIONAL_0_Z7771\: LUT5 
generic map(
  INIT => X"11111110"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS\,
  I1 => N_3812,
  I2 => \GRLFPC20.FPO.FRAC\(54),
  I3 => N_3881,
  I4 => N_3880,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN30_CONDITIONAL_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_SS0_Z7772\: LUT3 
generic map(
  INIT => X"CD"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST\(17),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST\(15),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_SS0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_SS9_Z7773\: LUT3 
generic map(
  INIT => X"BA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_3_REP1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_SS9\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1[0]_Z7774\: LUT5 
generic map(
  INIT => X"535CA3AC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
\GRLFPC20.COMB.DBGDATA_4[20]\: LUT4 
generic map(
  INIT => X"3210"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => rfo1_data1(20),
  I3 => rfo2_data1(20),
  O => cpo_dbg_data(20));
\GRLFPC20.COMB.DBGDATA_4[17]\: LUT4 
generic map(
  INIT => X"FEDC"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => rfo1_data1(17),
  I3 => rfo2_data1(17),
  O => cpo_dbg_data(17));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_21[75]\: LUT4_L 
generic map(
  INIT => X"A695"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(48),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(52),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8825\);
\GRLFPC20.COMB.DBGDATA_4[12]\: LUT4 
generic map(
  INIT => X"3210"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => rfo1_data1(12),
  I3 => rfo2_data1(12),
  O => cpo_dbg_data(12));
\GRLFPC20.COMB.DBGDATA_4[21]\: LUT4 
generic map(
  INIT => X"3210"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => rfo1_data1(21),
  I3 => rfo2_data1(21),
  O => cpo_dbg_data(21));
\GRLFPC20.COMB.DBGDATA_4[18]\: LUT4 
generic map(
  INIT => X"FEDC"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => rfo1_data1(18),
  I3 => rfo2_data1(18),
  O => cpo_dbg_data(18));
\GRLFPC20.COMB.DBGDATA_4[19]\: LUT4 
generic map(
  INIT => X"3210"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => rfo1_data1(19),
  I3 => rfo2_data1(19),
  O => cpo_dbg_data(19));
\GRLFPC20.COMB.DBGDATA_4[28]\: LUT4 
generic map(
  INIT => X"3210"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => rfo1_data1(28),
  I3 => rfo2_data1(28),
  O => cpo_dbg_data(28));
\GRLFPC20.COMB.DBGDATA_4[29]\: LUT4 
generic map(
  INIT => X"3210"
)
port map (
  I0 => cpi_dbg_addr(0),
  I1 => cpi_dbg_fsr,
  I2 => rfo1_data1(29),
  I3 => rfo2_data1(29),
  O => cpo_dbg_data(29));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4[3]_Z7784\: LUT5 
generic map(
  INIT => X"5A5A33CC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3[2]_Z7785\: LUT5 
generic map(
  INIT => X"53A35CAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2[1]_Z7786\: LUT5 
generic map(
  INIT => X"53A35CAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.UN198_TEMP_Z7787\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.UN198_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_1[5]\: LUT3_L 
generic map(
  INIT => X"80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRLOI\(30),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRLOI\(34),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRLOI\(29),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8537_RETI\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2[3]_Z7789\: LUT3 
generic map(
  INIT => X"CE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_30_REP1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_29_REP1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_FAST\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M8[2]_Z7790\: LUT3_L 
generic map(
  INIT => X"FE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_7_REP1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_8_REP1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_9_REP1\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M8\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD_Z7791\: LUT4 
generic map(
  INIT => X"ECA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST\(374),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(12),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(9),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(11),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\);
\GRLFPC20.WRADDR_0_SQMUXA_Z7792\: LUT3 
generic map(
  INIT => X"20"
)
port map (
  I0 => cpi_dbg_enable,
  I1 => cpi_dbg_fsr,
  I2 => cpi_dbg_write,
  O => \GRLFPC20.WRADDR_0_SQMUXA\);
\GRLFPC20.COMB.V.X.FPOP_1_Z7793\: LUT3_L 
generic map(
  INIT => X"10"
)
port map (
  I0 => cpi_m_annul,
  I1 => cpi_m_trap,
  I2 => \GRLFPC20.R.M.FPOP\,
  LO => \GRLFPC20.COMB.V.X.FPOP_1\);
\GRLFPC20.COMB.V.X.LD_1_Z7794\: LUT3_L 
generic map(
  INIT => X"10"
)
port map (
  I0 => cpi_m_annul,
  I1 => cpi_m_trap,
  I2 => \GRLFPC20.R.M.LD\,
  LO => \GRLFPC20.COMB.V.X.LD_1\);
\GRLFPC20.COMB.V.M.FPOP_1_Z7795\: LUT3_L 
generic map(
  INIT => X"10"
)
port map (
  I0 => cpi_e_annul,
  I1 => cpi_e_trap,
  I2 => \GRLFPC20.R.E.FPOP\,
  LO => \GRLFPC20.COMB.V.M.FPOP_1\);
\GRLFPC20.COMB.V.M.LD_1_Z7796\: LUT3_L 
generic map(
  INIT => X"10"
)
port map (
  I0 => cpi_e_annul,
  I1 => cpi_e_trap,
  I2 => \GRLFPC20.R.E.LD\,
  LO => \GRLFPC20.COMB.V.M.LD_1\);
\GRLFPC20.COMB.V.E.AFQ_1_Z7797\: LUT3_L 
generic map(
  INIT => X"10"
)
port map (
  I0 => cpi_a_annul,
  I1 => cpi_a_trap,
  I2 => \GRLFPC20.R.A.AFQ\,
  LO => \GRLFPC20.COMB.V.E.AFQ_1\);
\GRLFPC20.COMB.V.E.LD_1_Z7798\: LUT3_L 
generic map(
  INIT => X"10"
)
port map (
  I0 => cpi_a_annul,
  I1 => cpi_a_trap,
  I2 => \GRLFPC20.R.A.LD\,
  LO => \GRLFPC20.COMB.V.E.LD_1\);
\GRLFPC20.COMB.V.M.AFQ_1_Z7799\: LUT3_L 
generic map(
  INIT => X"10"
)
port map (
  I0 => cpi_e_annul,
  I1 => cpi_e_trap,
  I2 => \GRLFPC20.R.E.AFQ\,
  LO => \GRLFPC20.COMB.V.M.AFQ_1\);
\GRLFPC20.COMB.V.X.AFQ_1_Z7800\: LUT3_L 
generic map(
  INIT => X"10"
)
port map (
  I0 => cpi_m_annul,
  I1 => cpi_m_trap,
  I2 => \GRLFPC20.R.M.AFQ\,
  LO => \GRLFPC20.COMB.V.X.AFQ_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS_2[1]_Z7801\: LUT3 
generic map(
  INIT => X"E0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(3),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(5),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS_2\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0_0_A2_0_0[0]\: LUT4 
generic map(
  INIT => X"0004"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0_0_A2_0\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.REEXCOVUV.UN18_LOCOV_Z7803\: LUT3 
generic map(
  INIT => X"80"
)
port map (
  I0 => \GRLFPC20.FPO.EXP\(8),
  I1 => \GRLFPC20.FPO.EXP\(9),
  I2 => \GRLFPC20.FPO.EXP\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.REEXCOVUV.UN18_LOCOV\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.REEXCOVUV.UN25_LOCOV_Z7804\: LUT3 
generic map(
  INIT => X"FE"
)
port map (
  I0 => \GRLFPC20.FPO.EXP\(8),
  I1 => \GRLFPC20.FPO.EXP\(9),
  I2 => \GRLFPC20.FPO.EXP\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.REEXCOVUV.UN25_LOCOV\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_0_A2[1]\: LUT4_L 
generic map(
  INIT => X"0040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(41),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(38),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(39),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(40),
  LO => \GRLFPC20.FPO.EXC\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_0_A2[3]\: LUT3_L 
generic map(
  INIT => X"02"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(38),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(39),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(40),
  LO => \GRLFPC20.FPO.EXC\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_Z7807\: LUT4 
generic map(
  INIT => X"8000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(49),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(51),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(52),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(50),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_6_Z7808\: LUT4 
generic map(
  INIT => X"FFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_6\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_9_Z7809\: LUT4 
generic map(
  INIT => X"0001"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST\(3),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_9\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1_2[6]_Z7810\: LUT4_L 
generic map(
  INIT => X"FFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(254),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(253),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(255),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(256),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1_2\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN12_SRTOSTICKY_3_Z7811\: LUT4_L 
generic map(
  INIT => X"FFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(6),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(7),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(8),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(9),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN12_SRTOSTICKY_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_2_Z7812\: LUT3 
generic map(
  INIT => X"80"
)
port map (
  I0 => \GRLFPC20.FPO.FRAC\(50),
  I1 => \GRLFPC20.FPO.FRAC\(51),
  I2 => \GRLFPC20.FPO.FRAC\(54),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2[59]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(54),
  I2 => N_3881,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9127\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH[8]_Z7814\: LUT3 
generic map(
  INIT => X"E4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_FAST\(10),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2[58]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => N_3880,
  I2 => N_3882,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9128\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB[0]_Z7816\: LUT3 
generic map(
  INIT => X"D1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(19),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1[244]\: LUT3 
generic map(
  INIT => X"B8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(257),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
  I2 => \GRLFPC20.FPO.EXP\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8587\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2[63]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(50),
  I2 => \GRLFPC20.FPO.FRAC\(52),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9123\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2[61]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(52),
  I2 => \GRLFPC20.FPO.FRAC\(54),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9125\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIFJBB[69]\: LUT1_L 
generic map(
  INIT => X"1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(69),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(69));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_7_Z7821\: LUT2 
generic map(
  INIT => X"1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_7\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_2_2_0_O2[25]\: LUT2 
generic map(
  INIT => X"B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_746\);
\GRLFPC20.COMB.WREN12\: LUT2 
generic map(
  INIT => X"1"
)
port map (
  I0 => cpi_x_cnt(0),
  I1 => cpi_x_cnt(1),
  O => \GRLFPC20.N_2045\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SFTLFT.AREGXORBREG_Z7824\: LUT2_L 
generic map(
  INIT => X"6"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(13),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(12),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SFTLFT.AREGXORBREG\);
\GRLFPC20.R.I.EXC_RNIAG8C[4]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.R.I.EXC\(4),
  I1 => \GRLFPC20.R.FSR.TEM\(4),
  O => \GRLFPC20.N_1310\);
\GRLFPC20.R.I.EXC_RNI288C[0]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.R.I.EXC\(0),
  I1 => \GRLFPC20.R.FSR.TEM\(0),
  O => \GRLFPC20.N_1306\);
\GRLFPC20.R.I.EXC_RNI4A8C[1]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.R.I.EXC\(1),
  I1 => \GRLFPC20.R.FSR.TEM\(1),
  O => \GRLFPC20.N_1307\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_RNO[15]\: LUT1_L 
generic map(
  INIT => X"1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(42));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_12_Z7829\: LUT2 
generic map(
  INIT => X"9"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(232),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(245),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_12\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_RNO[11]\: LUT1_L 
generic map(
  INIT => X"1"
)
port map (
  I0 => cpi_d_inst(6),
  LO => CPI_D_INST_I(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.REEXCOVUV.UN13_LOCOV_0_2_Z7831\: LUT2_L 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.FPO.EXP\(5),
  I1 => \GRLFPC20.FPO.EXP\(6),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.REEXCOVUV.UN13_LOCOV_0_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0[58]_Z7832\: LUT6 
generic map(
  INIT => X"C0C0D5C0C0C0C0C0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A30_4_0\(58),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A30_4_1\(58),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9828\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12195\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10647\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0\(58));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNILCJQ1[62]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIVMJQ1[67]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI9JUM1[75]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI7J0N1[84]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIPKNQ1[83]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIUQOQ1[89]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI5J2N1[91]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.CIN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNISTKQ[110]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIN7BU[108]\: LUT5 
generic map(
  INIT => X"5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIV6SM1[62]\: LUT5 
generic map(
  INIT => X"3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5[52]_Z7843\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10211\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_715\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9454\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_1\(52),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4[6]_Z7844\: LUT6 
generic map(
  INIT => X"FFFFFFFF3B0A3300"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9506_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_143\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2708\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0\(6),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5[18]_Z7845\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF0040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9994_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_749\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1025\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0\(18),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5\(18));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7[53]_Z7846\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF08"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9503_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10236_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_906\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10299\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10294\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2\(53),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7\(53));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_11[57]_Z7847\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFF8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9975_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10626_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12238\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_1\(57),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_967\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2\(57),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_11\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"AC0053FF53FFAC00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.UN528_TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.UN531_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.SI_119\(50),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[51]\: LUT5 
generic map(
  INIT => X"3120FDEC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8313\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8315\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(52),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8636\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[13]\: LUT5 
generic map(
  INIT => X"3120FDEC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8351\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8353\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(14),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8674\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1_RNILJ132[33]\: LUT6 
generic map(
  INIT => X"7887788778788787"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\(33),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(33),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_33\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1_RNIMK132[34]\: LUT6 
generic map(
  INIT => X"7887788778788787"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\(34),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(34),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_34\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1_RNINL132[35]\: LUT6 
generic map(
  INIT => X"7887788778788787"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\(35),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(35),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_35\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1_RNI1V032[36]\: LUT6 
generic map(
  INIT => X"7887788778788787"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\(36),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(36),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_36\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1_RNI20132[37]\: LUT6 
generic map(
  INIT => X"7887788778788787"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\(37),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(37),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_37\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1_RNI31132[38]\: LUT6 
generic map(
  INIT => X"7887788778788787"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\(38),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(38),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_38\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1_RNIOO332[54]\: LUT6 
generic map(
  INIT => X"7887788778788787"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\(54),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(54),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_54\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1_LUT6_2_RNIUFE52[56]\: LUT6 
generic map(
  INIT => X"7887788778788787"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\(57),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(56),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_56\);
\GRLFPC20.RS1_1_0_0[3]_Z7859\: LUT5 
generic map(
  INIT => X"CAC0C0C0"
)
port map (
  I0 => cpi_d_inst(28),
  I1 => cpi_dbg_addr(3),
  I2 => cpi_dbg_enable,
  I3 => \GRLFPC20.RS1V_0_SQMUXA\,
  I4 => holdn,
  O => \GRLFPC20.RS1_1_0_0\(3));
\GRLFPC20.RS1_1_0_0[2]_Z7860\: LUT5 
generic map(
  INIT => X"CAC0C0C0"
)
port map (
  I0 => cpi_d_inst(27),
  I1 => cpi_dbg_addr(2),
  I2 => cpi_dbg_enable,
  I3 => \GRLFPC20.RS1V_0_SQMUXA\,
  I4 => holdn,
  O => \GRLFPC20.RS1_1_0_0\(2));
\GRLFPC20.RS1_1_0_0[1]_Z7861\: LUT5 
generic map(
  INIT => X"CAC0C0C0"
)
port map (
  I0 => cpi_d_inst(26),
  I1 => cpi_dbg_addr(1),
  I2 => cpi_dbg_enable,
  I3 => \GRLFPC20.RS1V_0_SQMUXA\,
  I4 => holdn,
  O => \GRLFPC20.RS1_1_0_0\(1));
\GRLFPC20.RS1_1_0_0[4]_Z7862\: LUT5 
generic map(
  INIT => X"CAC0C0C0"
)
port map (
  I0 => cpi_d_inst(29),
  I1 => cpi_dbg_addr(4),
  I2 => cpi_dbg_enable,
  I3 => \GRLFPC20.RS1V_0_SQMUXA\,
  I4 => holdn,
  O => \GRLFPC20.RS1_1_0_0\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[67]_Z7863\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(67),
    D => NN_4,
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_0_CY_Z7864\: MUXCY_L port map (
    DI => NN_2,
    CI => NN_3,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN8_TEMP\(0),
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_0_CY\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_0_CY_Z7865\: MUXCY_L port map (
    DI => NN_2,
    CI => NN_3,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.MIXOIN\(0),
    LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_0_CY\);
\GRLFPC20.V.I.V_3_SQMUXA_Z7866\: LUT6_L 
generic map(
  INIT => X"0000000000AA00A2"
)
port map (
  I0 => \GRLFPC20.V.I.V_3_SQMUXA_0\,
  I1 => \GRLFPC20.N_1837\,
  I2 => \GRLFPC20.COMB.V.STATE_9\(1),
  I3 => \GRLFPC20.COMB.ANNULRES_1\,
  I4 => \GRLFPC20.COMB.V.STATE_9\(0),
  I5 => \GRLFPC20.N_2112\,
  LO => \GRLFPC20.V.I.V_3_SQMUXA\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"9966966966996996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_AC0_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.SI_80\(33),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_AC0_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(24));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24.Z_C4\: LUT6 
generic map(
  INIT => X"EEBBEBBE88228228"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_AC0_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.SI_80\(33),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_AC0_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(81));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_19[0]_Z7869\: LUT5 
generic map(
  INIT => X"4D5F0517"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SBLSBS_1\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN16_NOTPROP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO1_0\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN18_GEN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_9\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_19\(0));
\GRLFPC20.COMB.V.MK.BUSY2_2_Z7870\: LUT6_L 
generic map(
  INIT => X"00000000084C0000"
)
port map (
  I0 => \GRLFPC20.N_1295\,
  I1 => \GRLFPC20.R.MK.BUSY\,
  I2 => \GRLFPC20.R.X.FPOP\,
  I3 => \GRLFPC20.R.X.SEQERR\,
  I4 => \GRLFPC20.N_1528\,
  I5 => \GRLFPC20.N_2015\,
  LO => \GRLFPC20.COMB.V.MK.BUSY2_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M_RNO[5]\: LUT5 
generic map(
  INIT => X"FFBF008F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14\(77),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN3_NOTRESETORUNIMP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8114\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_11\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_2\: LUT5 
generic map(
  INIT => X"0000A0A8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14_2\(77),
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14\(77),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_4_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.STKGEN_3_RNO\: LUT5 
generic map(
  INIT => X"DEED4884"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_453\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.SI_55\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_943_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1_RNISHHT6\: LUT6 
generic map(
  INIT => X"9669699669969669"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_453\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55.Z_C1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.SI_55\(2),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN22_NOTPROP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"399CC663C663399C"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_544\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.SI_44\(13),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44.Z_AXB2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(45));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45.Z_C4\: LUT6 
generic map(
  INIT => X"CEEFFDDC088CC440"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_544\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.SI_44\(13),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44.Z_AXB2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(102));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_1_A2_0_A2_LUT6_2_RNIAHJA3[56]\: LUT6 
generic map(
  INIT => X"0055000030753030"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_783\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_775\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2606\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_717\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2584\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1592\);
\GRLFPC20.R.A.FPOP_RNO\: LUT6_L 
generic map(
  INIT => X"0000000000000100"
)
port map (
  I0 => cpi_d_annul,
  I1 => cpi_d_trap,
  I2 => cpi_flush,
  I3 => \GRLFPC20.N_1583\,
  I4 => CPO_EXC_1,
  I5 => \GRLFPC20.COMB.LOCKGEN.LOCKI\,
  LO => \GRLFPC20.N_1312\);
\GRLFPC20.COMB.V.A.ST_1_Z7879\: LUT6_L 
generic map(
  INIT => X"0000000000000100"
)
port map (
  I0 => cpi_d_annul,
  I1 => cpi_d_trap,
  I2 => cpi_flush,
  I3 => \GRLFPC20.COMB.FPDECODE.ST\,
  I4 => CPO_EXC_1,
  I5 => \GRLFPC20.COMB.LOCKGEN.LOCKI\,
  LO => \GRLFPC20.COMB.V.A.ST_1\);
\GRLFPC20.COMB.V.A.AFQ_1_Z7880\: LUT6_L 
generic map(
  INIT => X"0000000000000100"
)
port map (
  I0 => cpi_d_annul,
  I1 => cpi_d_trap,
  I2 => cpi_flush,
  I3 => \GRLFPC20.COMB.V.A.AFQ_1_1\,
  I4 => CPO_EXC_1,
  I5 => \GRLFPC20.COMB.LOCKGEN.LOCKI\,
  LO => \GRLFPC20.COMB.V.A.AFQ_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[39]\: LUT5 
generic map(
  INIT => X"3120FDEC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8325\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8327\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(40),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8648\);
\GRLFPC20.R.A.RF2REN_RNO[1]\: LUT6_L 
generic map(
  INIT => X"00000000FFB80000"
)
port map (
  I0 => \GRLFPC20.COMB.FPDECODE.RS1D5\,
  I1 => \GRLFPC20.N_925\,
  I2 => \GRLFPC20.RS1D_CNST\,
  I3 => \GRLFPC20.N_2962\,
  I4 => \GRLFPC20.COMB.RS1V_1\,
  I5 => \GRLFPC20.COMB.LOCKGEN.LOCKI\,
  LO => \GRLFPC20.N_2961_I\);
\GRLFPC20.COMB.V.A.RF2REN_1[1]_Z7883\: LUT6 
generic map(
  INIT => X"0F0D00000F080000"
)
port map (
  I0 => \GRLFPC20.N_925\,
  I1 => \GRLFPC20.COMB.FPDECODE.RS1D5\,
  I2 => \GRLFPC20.COMB.LOCKGEN.LOCKI\,
  I3 => \GRLFPC20.COMB.RS1_1\(0),
  I4 => \GRLFPC20.COMB.RS1V_1\,
  I5 => \GRLFPC20.RS1D_CNST\,
  O => \GRLFPC20.COMB.V.A.RF2REN_1\(1));
\GRLFPC20.COMB.V.A.RF1REN_1[1]_Z7884\: LUT6 
generic map(
  INIT => X"0D0F0000080F0000"
)
port map (
  I0 => \GRLFPC20.N_925\,
  I1 => \GRLFPC20.COMB.FPDECODE.RS1D5\,
  I2 => \GRLFPC20.COMB.LOCKGEN.LOCKI\,
  I3 => \GRLFPC20.COMB.RS1_1\(0),
  I4 => \GRLFPC20.COMB.RS1V_1\,
  I5 => \GRLFPC20.RS1D_CNST\,
  O => \GRLFPC20.COMB.V.A.RF1REN_1\(1));
\GRLFPC20.WREN1_1_SQMUXA_Z7885\: LUT6 
generic map(
  INIT => X"0000000000200000"
)
port map (
  I0 => cpi_x_inst(20),
  I1 => \GRLFPC20.N_1295\,
  I2 => \GRLFPC20.N_1475\,
  I3 => \GRLFPC20.N_2015\,
  I4 => \GRLFPC20.N_2045\,
  I5 => \GRLFPC20.R.X.SEQERR\,
  O => \GRLFPC20.WREN1_1_SQMUXA\);
\GRLFPC20.COMB.WREN1_1_RNO\: LUT6 
generic map(
  INIT => X"0000000000000100"
)
port map (
  I0 => cpi_x_inst(20),
  I1 => cpi_x_inst(25),
  I2 => \GRLFPC20.N_1295\,
  I3 => \GRLFPC20.N_1475\,
  I4 => \GRLFPC20.N_2015\,
  I5 => \GRLFPC20.R.X.SEQERR\,
  O => \GRLFPC20.COMB.WREN1_2_M\);
\GRLFPC20.R.I.EXEC_RNO\: LUT6_L 
generic map(
  INIT => X"000000BF00000000"
)
port map (
  I0 => \GRLFPC20.N_1295\,
  I1 => \GRLFPC20.R.X.SEQERR\,
  I2 => \GRLFPC20.N_1494\,
  I3 => \GRLFPC20.COMB.V.I.EXEC_18_0_29_I_0\,
  I4 => \GRLFPC20.N_2015\,
  I5 => \GRLFPC20.COMB.V.FSR.AEXC_1_SN.N_7_MUX\,
  LO => \GRLFPC20.N_2929_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31.Z_C3_Z7888\: LUT5 
generic map(
  INIT => X"EDDE8448"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.SI_30\(27),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_C1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_28[75]\: LUT5_L 
generic map(
  INIT => X"FFFBF7F3"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(50),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CONDMUXMULXFF.UN5_NOTSQRTLFTCC\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14\(77),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8815\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8830\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12\(75));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33.Z_C4\: LUT6 
generic map(
  INIT => X"CDDFFEEC044CC880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.SI_32\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_AXB2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(90));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"366CC993C993366C"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.SI_32\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_AXB2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(33));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54.Z_AXBXC3\: LUT6 
generic map(
  INIT => X"6996966996696996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_AXB1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54.Z_C4\: LUT6 
generic map(
  INIT => X"BEEBEBBE28828228"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_AXB1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53.Z_C2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(111));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10.Z_AXBXC2\: LUT5 
generic map(
  INIT => X"96696996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.SI_9\(48),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.SI_125\(44));
\GRLFPC20.COMB.WRDATA_4[21]_Z7895\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(21),
  I3 => \GRLFPC20.R.I.RES\(50),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(21));
\GRLFPC20.COMB.WRDATA_4[57]_Z7896\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(54),
  I3 => \GRLFPC20.R.I.RES\(57),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(57));
\GRLFPC20.COMB.WRDATA_4[14]_Z7897\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(14),
  I3 => \GRLFPC20.R.I.RES\(43),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(14));
\GRLFPC20.COMB.WRDATA_4[13]_Z7898\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(13),
  I3 => \GRLFPC20.R.I.RES\(42),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(13));
\GRLFPC20.COMB.WRDATA_4[6]_Z7899\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(6),
  I3 => \GRLFPC20.R.I.RES\(35),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(6));
\GRLFPC20.COMB.WRDATA_4[60]_Z7900\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(57),
  I3 => \GRLFPC20.R.I.RES\(60),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(60));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_1[28]\: LUT6 
generic map(
  INIT => X"1100000011001000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2701\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_222\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2343\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0[56]\: LUT6 
generic map(
  INIT => X"FFFFFFF3FFFFFFF5"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8631\);
\GRLFPC20.COMB.WRDATA_4[7]_Z7903\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(7),
  I3 => \GRLFPC20.R.I.RES\(36),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(7));
\GRLFPC20.COMB.WRDATA_4[5]_Z7904\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(5),
  I3 => \GRLFPC20.R.I.RES\(34),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(5));
\GRLFPC20.COMB.WRDATA_4[2]_Z7905\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(2),
  I3 => \GRLFPC20.R.I.RES\(31),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(2));
\GRLFPC20.RS2_1[3]\: LUT6 
generic map(
  INIT => X"CAC0CAC0CFCFC0C0"
)
port map (
  I0 => cpi_d_inst(3),
  I1 => cpi_dbg_addr(3),
  I2 => cpi_dbg_enable,
  I3 => \GRLFPC20.N_1583\,
  I4 => \GRLFPC20.R.A.RS2\(3),
  I5 => holdn,
  O => RFI2_RD2ADDR_22);
\GRLFPC20.COMB.WRDATA_4[32]_Z7907\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(29),
  I3 => \GRLFPC20.R.I.RES\(32),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(32));
\GRLFPC20.COMB.WRDATA_4[24]_Z7908\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(24),
  I3 => \GRLFPC20.R.I.RES\(53),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(24));
\GRLFPC20.COMB.WRDATA_4[20]_Z7909\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(20),
  I3 => \GRLFPC20.R.I.RES\(49),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(20));
\GRLFPC20.COMB.WRDATA_4[19]_Z7910\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(19),
  I3 => \GRLFPC20.R.I.RES\(48),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[11]_Z7911\: LUT6 
generic map(
  INIT => X"000800FBFF08FFFB"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8300\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8353\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[33]_Z7912\: LUT6 
generic map(
  INIT => X"000800FBFF08FFFB"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8278\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8331\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(33));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[14]_Z7913\: LUT6 
generic map(
  INIT => X"0800FB0008FFFBFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8295\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8352\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(14));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[15]_Z7914\: LUT6 
generic map(
  INIT => X"0800FB0008FFFBFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8294\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8351\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(15));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[38]_Z7915\: LUT6 
generic map(
  INIT => X"000800FBFF08FFFB"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8273\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8326\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(38));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[40]_Z7916\: LUT6 
generic map(
  INIT => X"0800FB0008FFFBFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8269\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8326\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(40));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[42]_Z7917\: LUT6 
generic map(
  INIT => X"000800FBFF08FFFB"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8269\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8322\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(42));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26[34]_Z7918\: LUT6 
generic map(
  INIT => X"0800FB0008FFFBFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8275\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8332\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(34));
\GRLFPC20.COMB.WRDATA_4[17]_Z7919\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(17),
  I3 => \GRLFPC20.R.I.RES\(46),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(17));
\GRLFPC20.COMB.WRDATA_4[16]_Z7920\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(16),
  I3 => \GRLFPC20.R.I.RES\(45),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(16));
\GRLFPC20.COMB.WRDATA_4[12]_Z7921\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(12),
  I3 => \GRLFPC20.R.I.RES\(41),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(12));
\GRLFPC20.COMB.WRDATA_4[54]_Z7922\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(51),
  I3 => \GRLFPC20.R.I.RES\(54),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(54));
\GRLFPC20.COMB.WRDATA_4[28]_Z7923\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(28),
  I3 => \GRLFPC20.R.I.RES\(57),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(28));
\GRLFPC20.COMB.WRDATA_4[26]_Z7924\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(26),
  I3 => \GRLFPC20.R.I.RES\(55),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(26));
\GRLFPC20.COMB.WRDATA_4[18]_Z7925\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(18),
  I3 => \GRLFPC20.R.I.RES\(47),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(18));
\GRLFPC20.COMB.WRDATA_4[15]_Z7926\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(15),
  I3 => \GRLFPC20.R.I.RES\(44),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(15));
\GRLFPC20.COMB.WRDATA_4[9]_Z7927\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(9),
  I3 => \GRLFPC20.R.I.RES\(38),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(9));
\GRLFPC20.COMB.WRDATA_4[4]_Z7928\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(4),
  I3 => \GRLFPC20.R.I.RES\(33),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(4));
\GRLFPC20.COMB.WRDATA_4[3]_Z7929\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(3),
  I3 => \GRLFPC20.R.I.RES\(32),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(3));
\GRLFPC20.COMB.WRDATA_4[1]_Z7930\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(1),
  I3 => \GRLFPC20.R.I.RES\(30),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(1));
\GRLFPC20.COMB.WRDATA_4[31]_Z7931\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(31),
  I3 => \GRLFPC20.R.I.RES\(63),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(31));
\GRLFPC20.RS2_1[1]\: LUT6 
generic map(
  INIT => X"CAC0CAC0CFCFC0C0"
)
port map (
  I0 => cpi_d_inst(1),
  I1 => cpi_dbg_addr(1),
  I2 => cpi_dbg_enable,
  I3 => \GRLFPC20.N_1583\,
  I4 => \GRLFPC20.R.A.RS2\(1),
  I5 => holdn,
  O => RFI2_RD2ADDR_20);
\GRLFPC20.COMB.WRDATA_4[8]_Z7933\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(8),
  I3 => \GRLFPC20.R.I.RES\(37),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(8));
\GRLFPC20.COMB.WRDATA_4[44]_Z7934\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(41),
  I3 => \GRLFPC20.R.I.RES\(44),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(44));
\GRLFPC20.COMB.WRDATA_4[25]_Z7935\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(25),
  I3 => \GRLFPC20.R.I.RES\(54),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(25));
\GRLFPC20.COMB.WRDATA_4[23]_Z7936\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(23),
  I3 => \GRLFPC20.R.I.RES\(52),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(23));
\GRLFPC20.COMB.WRDATA_4[22]_Z7937\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(22),
  I3 => \GRLFPC20.R.I.RES\(51),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(22));
\GRLFPC20.COMB.WRDATA_4[61]_Z7938\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(58),
  I3 => \GRLFPC20.R.I.RES\(61),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(61));
\GRLFPC20.COMB.WRDATA_4[59]_Z7939\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(56),
  I3 => \GRLFPC20.R.I.RES\(59),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(59));
\GRLFPC20.COMB.WRDATA_4[55]_Z7940\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(52),
  I3 => \GRLFPC20.R.I.RES\(55),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(55));
\GRLFPC20.COMB.WRDATA_4[0]_Z7941\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(0),
  I3 => \GRLFPC20.R.I.RES\(29),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(0));
\GRLFPC20.COMB.WRDATA_4[30]_Z7942\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(30),
  I3 => \GRLFPC20.R.I.RES\(59),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(30));
\GRLFPC20.RS2_1[2]\: LUT6 
generic map(
  INIT => X"CAC0CAC0CFCFC0C0"
)
port map (
  I0 => cpi_d_inst(2),
  I1 => cpi_dbg_addr(2),
  I2 => cpi_dbg_enable,
  I3 => \GRLFPC20.N_1583\,
  I4 => \GRLFPC20.R.A.RS2\(2),
  I5 => holdn,
  O => RFI2_RD2ADDR_21);
\GRLFPC20.COMB.WRDATA_4[10]_Z7944\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(10),
  I3 => \GRLFPC20.R.I.RES\(39),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(10));
\GRLFPC20.COMB.WRDATA_4[53]_Z7945\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(50),
  I3 => \GRLFPC20.R.I.RES\(53),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(53));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_AXB2_Z7946\: LUT6 
generic map(
  INIT => X"9669699669969669"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(21),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(21),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.CIN_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_552\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42.Z_AXB2\);
\GRLFPC20.RS2_1[4]\: LUT6 
generic map(
  INIT => X"CAC0CAC0CFCFC0C0"
)
port map (
  I0 => cpi_d_inst(4),
  I1 => cpi_dbg_addr(4),
  I2 => cpi_dbg_enable,
  I3 => \GRLFPC20.N_1583\,
  I4 => \GRLFPC20.R.A.RS2\(4),
  I5 => holdn,
  O => RFI2_RD2ADDR_23);
\GRLFPC20.COMB.WRDATA_4[39]_Z7948\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(36),
  I3 => \GRLFPC20.R.I.RES\(39),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(39));
\GRLFPC20.COMB.WRDATA_4[56]_Z7949\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(53),
  I3 => \GRLFPC20.R.I.RES\(56),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(56));
\GRLFPC20.COMB.WRDATA_4[62]_Z7950\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(59),
  I3 => \GRLFPC20.R.I.RES\(62),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(62));
\GRLFPC20.COMB.WRDATA_4[58]_Z7951\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(55),
  I3 => \GRLFPC20.R.I.RES\(58),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(58));
\GRLFPC20.COMB.WRDATA_4[11]_Z7952\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(11),
  I3 => \GRLFPC20.R.I.RES\(40),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(11));
\GRLFPC20.COMB.WRDATA_4[42]_Z7953\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(39),
  I3 => \GRLFPC20.R.I.RES\(42),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(42));
\GRLFPC20.COMB.WRDATA_4[41]_Z7954\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(38),
  I3 => \GRLFPC20.R.I.RES\(41),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(41));
\GRLFPC20.COMB.WRDATA_4[51]_Z7955\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(48),
  I3 => \GRLFPC20.R.I.RES\(51),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(51));
\GRLFPC20.COMB.WRDATA_4[49]_Z7956\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(46),
  I3 => \GRLFPC20.R.I.RES\(49),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(49));
\GRLFPC20.COMB.WRDATA_4[48]_Z7957\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(45),
  I3 => \GRLFPC20.R.I.RES\(48),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(48));
\GRLFPC20.COMB.WRDATA_4[45]_Z7958\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(42),
  I3 => \GRLFPC20.R.I.RES\(45),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(45));
\GRLFPC20.COMB.WRDATA_4[46]_Z7959\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(43),
  I3 => \GRLFPC20.R.I.RES\(46),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(46));
\GRLFPC20.COMB.WRDATA_4[43]_Z7960\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(40),
  I3 => \GRLFPC20.R.I.RES\(43),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(43));
\GRLFPC20.COMB.WRDATA_4[37]_Z7961\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(34),
  I3 => \GRLFPC20.R.I.RES\(37),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(37));
\GRLFPC20.COMB.WRDATA_4[36]_Z7962\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(33),
  I3 => \GRLFPC20.R.I.RES\(36),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(36));
\GRLFPC20.COMB.WRDATA_4[34]_Z7963\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(31),
  I3 => \GRLFPC20.R.I.RES\(34),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(34));
\GRLFPC20.COMB.WRDATA_4[33]_Z7964\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(30),
  I3 => \GRLFPC20.R.I.RES\(33),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(33));
\GRLFPC20.COMB.WRDATA_4[29]_Z7965\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(29),
  I3 => \GRLFPC20.R.I.RES\(58),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(29));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_2[50]\: LUT6 
generic map(
  INIT => X"0000802000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1232\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2151\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6.Z_AXB2_Z7967\: LUT6 
generic map(
  INIT => X"6996966996696996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(57),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.CIN_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6.Z_AXB2\);
\GRLFPC20.COMB.WRDATA_4[47]_Z7968\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(44),
  I3 => \GRLFPC20.R.I.RES\(47),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIJKU72[66]\: LUT6 
generic map(
  INIT => X"00000000FFFFFAF2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(66),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(67),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.ENTRYPOINT\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14\(77),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_0_SN_N_7_MUX\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38.Z_C2_Z7970\: LUT6 
generic map(
  INIT => X"FF2DFFD22D00D200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(349),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(24),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.CIN_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.CIN_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31.Z_C2_Z7971\: LUT6 
generic map(
  INIT => X"FF2DFFD22D00D200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(342),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(31),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.CIN_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.CIN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31.Z_C2\);
\GRLFPC20.COMB.WRDATA_4[27]_Z7972\: LUT6 
generic map(
  INIT => X"F1E0FB40F3C0F3C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(27),
  I3 => \GRLFPC20.R.I.RES\(56),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(27));
\GRLFPC20.COMB.WRDATA_4[40]_Z7973\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(37),
  I3 => \GRLFPC20.R.I.RES\(40),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(40));
\GRLFPC20.COMB.WRDATA_4[50]_Z7974\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(47),
  I3 => \GRLFPC20.R.I.RES\(50),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(50));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_12[29]\: LUT5 
generic map(
  INIT => X"00002000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_742\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2335\);
\GRLFPC20.COMB.WRDATA_4[35]_Z7976\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(32),
  I3 => \GRLFPC20.R.I.RES\(35),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(35));
\GRLFPC20.COMB.WRDATA_4[38]_Z7977\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(35),
  I3 => \GRLFPC20.R.I.RES\(38),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(38));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_RNO[12]\: LUT6 
generic map(
  INIT => X"0000000020000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_742\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_965\);
\GRLFPC20.COMB.WRDATA_4[52]_Z7979\: LUT6 
generic map(
  INIT => X"FE10F4B0FC30FC30"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.I.V\,
  I1 => \GRLFPC20.R.I.RDD\,
  I2 => \GRLFPC20.R.I.RES\(49),
  I3 => \GRLFPC20.R.I.RES\(52),
  I4 => \GRLFPC20.R.X.RDD\,
  I5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
  O => \GRLFPC20.COMB.WRDATA_4\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19[68]_Z7980\: LUT6 
generic map(
  INIT => X"FF00F0F0CCCCAAAA"
)
port map (
  I0 => rfo1_data1(12),
  I1 => rfo1_data1(15),
  I2 => rfo2_data1(12),
  I3 => rfo2_data1(15),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I5 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(68));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19[63]_Z7981\: LUT6 
generic map(
  INIT => X"FF00F0F0CCCCAAAA"
)
port map (
  I0 => rfo1_data1(17),
  I1 => rfo1_data1(20),
  I2 => rfo2_data1(17),
  I3 => rfo2_data1(20),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I5 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(63));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19[65]_Z7982\: LUT6 
generic map(
  INIT => X"FF00F0F0CCCCAAAA"
)
port map (
  I0 => rfo1_data1(15),
  I1 => rfo1_data1(18),
  I2 => rfo2_data1(15),
  I3 => rfo2_data1(18),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I5 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(65));
\GRLFPC20.COMB.V.E.STDATA_1_1[4]\: LUT5_L 
generic map(
  INIT => X"F0CCF0AA"
)
port map (
  I0 => rfo1_data1(4),
  I1 => rfo2_data1(4),
  I2 => \GRLFPC20.R.FSR.CEXC\(4),
  I3 => \GRLFPC20.R.A.AFSR\,
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  LO => \GRLFPC20.N_2376\);
\GRLFPC20.COMB.V.E.STDATA_1_1[30]\: LUT5_L 
generic map(
  INIT => X"F0CCF0AA"
)
port map (
  I0 => rfo1_data1(30),
  I1 => rfo2_data1(30),
  I2 => \GRLFPC20.R.FSR.RD\(0),
  I3 => \GRLFPC20.R.A.AFSR\,
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  LO => \GRLFPC20.N_2402\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19[82]_Z7985\: LUT5 
generic map(
  INIT => X"CCF0AAF0"
)
port map (
  I0 => rfo1_data1(1),
  I1 => rfo2_data1(1),
  I2 => rfo2_data1(30),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(82));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_1_1[32]_Z7986\: LUT6_L 
generic map(
  INIT => X"000000004000C000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_717\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_1_1\(32));
\GRLFPC20.COMB.RDD_2_Z7987\: LUT6 
generic map(
  INIT => X"F1F0F0F0E0F0F0F0"
)
port map (
  I0 => \GRLFPC20.N_1295\,
  I1 => \GRLFPC20.R.I.EXEC\,
  I2 => \GRLFPC20.R.I.RDD\,
  I3 => \GRLFPC20.R.I.V\,
  I4 => \GRLFPC20.R.X.FPOP\,
  I5 => \GRLFPC20.R.X.RDD\,
  O => \GRLFPC20.COMB.RDD_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51.Z_AC0_2_Z7988\: LUT6 
generic map(
  INIT => X"CC5A000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_812_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.SI_51\(6),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51.Z_AC0_2\);
\GRLFPC20.COMB.RDD_1.M4_E_I_A3_1_0\: LUT6 
generic map(
  INIT => X"0200000000000000"
)
port map (
  I0 => cpi_d_inst(5),
  I1 => cpi_d_inst(6),
  I2 => cpi_d_inst(7),
  I3 => cpi_d_inst(8),
  I4 => cpi_d_inst(11),
  I5 => \GRLFPC20.N_3116\,
  O => \GRLFPC20.N_3082\);
\GRLFPC20.COMB.V.A.RF2REN_1[2]_Z7990\: LUT6 
generic map(
  INIT => X"0F080F080F0F0F00"
)
port map (
  I0 => cpi_d_inst(0),
  I1 => \GRLFPC20.N_1583\,
  I2 => \GRLFPC20.COMB.LOCKGEN.LOCKI\,
  I3 => \GRLFPC20.COMB.RS2D_1\,
  I4 => \GRLFPC20.R.A.RS2\(0),
  I5 => holdn,
  O => \GRLFPC20.COMB.V.A.RF2REN_1\(2));
\GRLFPC20.COMB.V.A.RF1REN_1DUP[2]\: LUT6 
generic map(
  INIT => X"0C040C040C000C0C"
)
port map (
  I0 => cpi_d_inst(0),
  I1 => \GRLFPC20.N_1583\,
  I2 => \GRLFPC20.COMB.LOCKGEN.LOCKI\,
  I3 => \GRLFPC20.COMB.RS2D_1\,
  I4 => \GRLFPC20.R.A.RS2\(0),
  I5 => holdn,
  O => N_11445);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19[61]_Z7992\: LUT6 
generic map(
  INIT => X"FF00F0F0CCCCAAAA"
)
port map (
  I0 => rfo1_data1(19),
  I1 => rfo1_data1(22),
  I2 => rfo2_data1(19),
  I3 => rfo2_data1(22),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I5 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(61));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_RNO[18]\: LUT6 
generic map(
  INIT => X"B1F0000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10207_I_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9858_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1036\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_12[13]\: LUT6 
generic map(
  INIT => X"0020000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10025_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9561\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_AC0_2_Z7995\: LUT6 
generic map(
  INIT => X"CC5A000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_846_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.SI_25\(32),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_AC0_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIA8B14[78]\: LUT6 
generic map(
  INIT => X"0000000000000010"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10410\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_966\);
\GRLFPC20.COMB.FPDECODE.RS1D5_0_A3\: LUT6 
generic map(
  INIT => X"0004000000000000"
)
port map (
  I0 => cpi_d_inst(8),
  I1 => cpi_d_inst(9),
  I2 => cpi_d_inst(12),
  I3 => cpi_d_inst(13),
  I4 => \GRLFPC20.N_3117\,
  I5 => \GRLFPC20.N_3120\,
  O => \GRLFPC20.COMB.FPDECODE.RS1D5\);
\GRLFPC20.COMB.RS1_1[0]_Z7998\: LUT6 
generic map(
  INIT => X"AFAFCF0FA0A0C000"
)
port map (
  I0 => cpi_d_inst(14),
  I1 => cpi_d_inst(25),
  I2 => holdn,
  I3 => \GRLFPC20.RS1V_0_SQMUXA\,
  I4 => \GRLFPC20.N_1583\,
  I5 => \GRLFPC20.R.A.RS1\(0),
  O => \GRLFPC20.COMB.RS1_1\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_20[6]\: LUT6 
generic map(
  INIT => X"0000000800000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9972_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9511\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15[2]\: LUT6 
generic map(
  INIT => X"0600000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9506_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9861_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2565\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A14_3[34]\: LUT6_L 
generic map(
  INIT => X"0000400000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9601_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9968\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_A26_23[31]\: LUT6 
generic map(
  INIT => X"0000000000000080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9409\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19[83]_Z8003\: LUT5 
generic map(
  INIT => X"CCF0AAF0"
)
port map (
  I0 => rfo1_data1(0),
  I1 => rfo2_data1(0),
  I2 => rfo2_data1(29),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I4 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(83));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A12_8[0]\: LUT6 
generic map(
  INIT => X"0200000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_314_I\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9454\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2[44]\: LUT6 
generic map(
  INIT => X"0000000000000040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_715\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2734\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_18[55]\: LUT6 
generic map(
  INIT => X"4000000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9655_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10456\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_13[32]\: LUT6 
generic map(
  INIT => X"0000000002000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10410\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9860\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A24_4[59]\: LUT6 
generic map(
  INIT => X"0000000022030000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9610_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_406\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10751\);
\GRLFPC20.COMB.V.FSR.AEXC_1_M0[2]_Z8009\: LUT5 
generic map(
  INIT => X"E2F0F0F0"
)
port map (
  I0 => cpi_lddata(7),
  I1 => \GRLFPC20.N_1295\,
  I2 => \GRLFPC20.R.FSR.AEXC\(2),
  I3 => \GRLFPC20.R.X.AFSR\,
  I4 => \GRLFPC20.R.X.LD\,
  O => \GRLFPC20.COMB.V.FSR.AEXC_1_M0\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_23[11]\: LUT6 
generic map(
  INIT => X"0000000000000008"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9666_1_I_0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9338\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_20[55]\: LUT6 
generic map(
  INIT => X"0008000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10888_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10458\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_15[13]\: LUT6 
generic map(
  INIT => X"0010000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9610_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12249\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_7_0_A2[49]\: LUT6 
generic map(
  INIT => X"0000000800000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2166\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_0_0_A2[16]\: LUT6 
generic map(
  INIT => X"00000000000B0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_291_I\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9666_1_I_0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_534\);
\GRLFPC20.COMB.V.FSR.AEXC_1_M0[4]_Z8015\: LUT5 
generic map(
  INIT => X"E2F0F0F0"
)
port map (
  I0 => cpi_lddata(9),
  I1 => \GRLFPC20.N_1295\,
  I2 => \GRLFPC20.R.FSR.AEXC\(4),
  I3 => \GRLFPC20.R.X.AFSR\,
  I4 => \GRLFPC20.R.X.LD\,
  O => \GRLFPC20.COMB.V.FSR.AEXC_1_M0\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_3[6]\: LUT6_L 
generic map(
  INIT => X"1000100000001000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9494\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19[79]_Z8017\: LUT6 
generic map(
  INIT => X"FF00F0F0CCCCAAAA"
)
port map (
  I0 => rfo1_data1(1),
  I1 => rfo1_data1(4),
  I2 => rfo2_data1(1),
  I3 => rfo2_data1(4),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I5 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(79));
\GRLFPC20.COMB.V.FSR.AEXC_1_M0[3]_Z8018\: LUT5 
generic map(
  INIT => X"E2F0F0F0"
)
port map (
  I0 => cpi_lddata(8),
  I1 => \GRLFPC20.N_1295\,
  I2 => \GRLFPC20.R.FSR.AEXC\(3),
  I3 => \GRLFPC20.R.X.AFSR\,
  I4 => \GRLFPC20.R.X.LD\,
  O => \GRLFPC20.COMB.V.FSR.AEXC_1_M0\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A26_8[60]\: LUT6_L 
generic map(
  INIT => X"0000000011010000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10827\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_0[49]\: LUT6 
generic map(
  INIT => X"0000000012001300"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_717\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2159\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_12[24]\: LUT6 
generic map(
  INIT => X"00200000002000A0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1187\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_1[36]\: LUT6_L 
generic map(
  INIT => X"D202000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9738_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10023\);
\GRLFPC20.COMB.V.FSR.AEXC_1_M0[0]_Z8023\: LUT5 
generic map(
  INIT => X"E2F0F0F0"
)
port map (
  I0 => cpi_lddata(5),
  I1 => \GRLFPC20.N_1295\,
  I2 => \GRLFPC20.R.FSR.AEXC\(0),
  I3 => \GRLFPC20.R.X.AFSR\,
  I4 => \GRLFPC20.R.X.LD\,
  O => \GRLFPC20.COMB.V.FSR.AEXC_1_M0\(0));
\GRLFPC20.COMB.V.FSR.FCC_1_M0[1]_Z8024\: LUT5 
generic map(
  INIT => X"E2F0F0F0"
)
port map (
  I0 => cpi_lddata(11),
  I1 => \GRLFPC20.N_1295\,
  I2 => CPO_CC_3,
  I3 => \GRLFPC20.R.X.AFSR\,
  I4 => \GRLFPC20.R.X.LD\,
  O => \GRLFPC20.COMB.V.FSR.FCC_1_M0\(1));
\GRLFPC20.COMB.V.FSR.FCC_1_M0[0]_Z8025\: LUT5 
generic map(
  INIT => X"E2F0F0F0"
)
port map (
  I0 => cpi_lddata(10),
  I1 => \GRLFPC20.N_1295\,
  I2 => NN_1,
  I3 => \GRLFPC20.R.X.AFSR\,
  I4 => \GRLFPC20.R.X.LD\,
  O => \GRLFPC20.COMB.V.FSR.FCC_1_M0\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_24[33]\: LUT6 
generic map(
  INIT => X"0000000000800000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9506_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10410\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9928\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_7[50]\: LUT6 
generic map(
  INIT => X"0000000000008000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2156\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_10[61]\: LUT6 
generic map(
  INIT => X"0000000000200000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9558_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_720\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10893\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_A2[20]\: LUT6 
generic map(
  INIT => X"0000000000002080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_717\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_720\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1034\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A22_19[53]\: LUT6 
generic map(
  INIT => X"0002000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9667_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9600_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10310\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_17[58]\: LUT6 
generic map(
  INIT => X"0000000020000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9558_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1971\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15[38]\: LUT6 
generic map(
  INIT => X"0000000000008200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_409\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10410\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2235\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_0[29]\: LUT6 
generic map(
  INIT => X"0000000000000040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10410\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2336\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_A2_2[37]\: LUT6 
generic map(
  INIT => X"0000000000004000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_749\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_720\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_972\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_0_A2_0_A2[40]\: LUT6 
generic map(
  INIT => X"0000000000002000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10410\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2230\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A22_13[53]\: LUT6 
generic map(
  INIT => X"0400000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10304\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A22_14[53]\: LUT6 
generic map(
  INIT => X"0000000040000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10305\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_8_3[36]\: LUT4 
generic map(
  INIT => X"8000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10030_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A26_15[56]\: LUT6 
generic map(
  INIT => X"2220000000200000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10535\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A26_5[60]\: LUT6 
generic map(
  INIT => X"2112000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10824\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.UN636_TEMP_Z8041\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.UN636_TEMP\);
\GRLFPC20.FPI.OP1[52]_Z8042\: LUT6 
generic map(
  INIT => X"E4E4F0CCCCCCF0CC"
)
port map (
  I0 => cpi_a_cnt(1),
  I1 => rfo1_data1(20),
  I2 => rfo2_data1(20),
  I3 => \GRLFPC20.R.A.RS1\(0),
  I4 => \GRLFPC20.R.A.RS1D\,
  I5 => \GRLFPC20.R.A.ST\,
  O => \GRLFPC20.FPI.OP1\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI0P1B1[99]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(16));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI02QS[101]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(14));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIRJ1B1[94]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(21));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A22_2_0[53]_Z8046\: LUT5_L 
generic map(
  INIT => X"00A000C0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A22_2_0\(53));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_10_A2_0_A2[60]\: LUT4 
generic map(
  INIT => X"1000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2602\);
\GRLFPC20.FPI.OP1[62]_Z8048\: LUT6 
generic map(
  INIT => X"E4E4F0CCCCCCF0CC"
)
port map (
  I0 => cpi_a_cnt(1),
  I1 => rfo1_data1(30),
  I2 => rfo2_data1(30),
  I3 => \GRLFPC20.R.A.RS1\(0),
  I4 => \GRLFPC20.R.A.RS1D\,
  I5 => \GRLFPC20.R.A.ST\,
  O => \GRLFPC20.FPI.OP1\(62));
\GRLFPC20.FPI.OP1[53]_Z8049\: LUT6 
generic map(
  INIT => X"E4E4F0CCCCCCF0CC"
)
port map (
  I0 => cpi_a_cnt(1),
  I1 => rfo1_data1(21),
  I2 => rfo2_data1(21),
  I3 => \GRLFPC20.R.A.RS1\(0),
  I4 => \GRLFPC20.R.A.RS1D\,
  I5 => \GRLFPC20.R.A.ST\,
  O => \GRLFPC20.FPI.OP1\(53));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIUL0B1[88]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(27));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0[236]_Z8051\: LUT6 
generic map(
  INIT => X"00CC00AAF0F0F0F0"
)
port map (
  I0 => rfo1_data2(28),
  I1 => rfo2_data2(28),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(236),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I4 => \GRLFPC20.COMB.UN1_FPCI_4\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8580\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_8_1[19]_Z8052\: LUT5 
generic map(
  INIT => X"03000100"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_8_1\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_1_1[7]_Z8053\: LUT6 
generic map(
  INIT => X"0000000000004080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_1_1\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNISK1B1[95]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(20));
\GRLFPC20.COMB.V.E.STDATA_1_0[15]\: LUT4 
generic map(
  INIT => X"F2D0"
)
port map (
  I0 => cpi_a_cnt(0),
  I1 => cpi_a_cnt(1),
  I2 => \GRLFPC20.R.I.INST\(15),
  I3 => \GRLFPC20.R.I.PC\(15),
  O => \GRLFPC20.N_2354\);
\GRLFPC20.COMB.V.E.STDATA_1_0[8]\: LUT4 
generic map(
  INIT => X"F2D0"
)
port map (
  I0 => cpi_a_cnt(0),
  I1 => cpi_a_cnt(1),
  I2 => \GRLFPC20.R.I.INST\(8),
  I3 => \GRLFPC20.R.I.PC\(8),
  O => \GRLFPC20.N_2347\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A30_10_1[58]_Z8057\: LUT5_L 
generic map(
  INIT => X"20000200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A30_10_1\(58));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_0[56]_Z8058\: LUT6 
generic map(
  INIT => X"C300C20000000002"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_0\(56));
\GRLFPC20.FPI.OP1[60]_Z8059\: LUT6 
generic map(
  INIT => X"E4E4F0CCCCCCF0CC"
)
port map (
  I0 => cpi_a_cnt(1),
  I1 => rfo1_data1(28),
  I2 => rfo2_data1(28),
  I3 => \GRLFPC20.R.A.RS1\(0),
  I4 => \GRLFPC20.R.A.RS1D\,
  I5 => \GRLFPC20.R.A.ST\,
  O => \GRLFPC20.FPI.OP1\(60));
\GRLFPC20.FPI.OP1[49]_Z8060\: LUT6 
generic map(
  INIT => X"E4E4F0CCCCCCF0CC"
)
port map (
  I0 => cpi_a_cnt(1),
  I1 => rfo1_data1(17),
  I2 => rfo2_data1(17),
  I3 => \GRLFPC20.R.A.RS1\(0),
  I4 => \GRLFPC20.R.A.RS1D\,
  I5 => \GRLFPC20.R.A.ST\,
  O => \GRLFPC20.FPI.OP1\(49));
\GRLFPC20.FPI.OP1[44]_Z8061\: LUT6 
generic map(
  INIT => X"E4E4F0CCCCCCF0CC"
)
port map (
  I0 => cpi_a_cnt(1),
  I1 => rfo1_data1(12),
  I2 => rfo2_data1(12),
  I3 => \GRLFPC20.R.A.RS1\(0),
  I4 => \GRLFPC20.R.A.RS1D\,
  I5 => \GRLFPC20.R.A.ST\,
  O => \GRLFPC20.FPI.OP1\(44));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0[234]_Z8062\: LUT6 
generic map(
  INIT => X"00CC00AAF0F0F0F0"
)
port map (
  I0 => rfo1_data2(30),
  I1 => rfo2_data2(30),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(234),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I4 => \GRLFPC20.COMB.UN1_FPCI_4\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8582\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_1[29]\: LUT6 
generic map(
  INIT => X"0000020000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2818\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_I_18\: LUT6 
generic map(
  INIT => X"A695596A00000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8554\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8539\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(9),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_I_18_0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_N_18\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_8_1[13]_Z8065\: LUT5 
generic map(
  INIT => X"04000100"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_8_1\(13));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIPK4R[246]\: LUT4 
generic map(
  INIT => X"C0A0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(233),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(246),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_I_5\: LUT5_L 
generic map(
  INIT => X"A695596A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8546\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8533\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12041\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI76MH1[255]\: LUT6 
generic map(
  INIT => X"AAAAFFF0CCCC0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(255),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(242),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(2));
\GRLFPC20.FPI.OP1[61]_Z8069\: LUT6 
generic map(
  INIT => X"E4E4F0CCCCCCF0CC"
)
port map (
  I0 => cpi_a_cnt(1),
  I1 => rfo1_data1(29),
  I2 => rfo2_data1(29),
  I3 => \GRLFPC20.R.A.RS1\(0),
  I4 => \GRLFPC20.R.A.RS1D\,
  I5 => \GRLFPC20.R.A.ST\,
  O => \GRLFPC20.FPI.OP1\(61));
\GRLFPC20.FPI.OP1[54]_Z8070\: LUT6 
generic map(
  INIT => X"E4E4F0CCCCCCF0CC"
)
port map (
  I0 => cpi_a_cnt(1),
  I1 => rfo1_data1(22),
  I2 => rfo2_data1(22),
  I3 => \GRLFPC20.R.A.RS1\(0),
  I4 => \GRLFPC20.R.A.RS1D\,
  I5 => \GRLFPC20.R.A.ST\,
  O => \GRLFPC20.FPI.OP1\(54));
\GRLFPC20.FPI.OP1[50]_Z8071\: LUT6 
generic map(
  INIT => X"E4E4F0CCCCCCF0CC"
)
port map (
  I0 => cpi_a_cnt(1),
  I1 => rfo1_data1(18),
  I2 => rfo2_data1(18),
  I3 => \GRLFPC20.R.A.RS1\(0),
  I4 => \GRLFPC20.R.A.RS1D\,
  I5 => \GRLFPC20.R.A.ST\,
  O => \GRLFPC20.FPI.OP1\(50));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIUM1B1[97]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(18));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNITL1B1[96]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNINF1B1[90]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(25));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIVM0B1[89]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(26));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_RNINE0B1[4]\: LUT4 
generic map(
  INIT => X"CCA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(4),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(31));
\GRLFPC20.FPI.OP1[38]_Z8077\: LUT6 
generic map(
  INIT => X"E4E4F0CCCCCCF0CC"
)
port map (
  I0 => cpi_a_cnt(1),
  I1 => rfo1_data1(6),
  I2 => rfo2_data1(6),
  I3 => \GRLFPC20.R.A.RS1\(0),
  I4 => \GRLFPC20.R.A.RS1D\,
  I5 => \GRLFPC20.R.A.ST\,
  O => \GRLFPC20.FPI.OP1\(38));
\GRLFPC20.FPI.OP1[40]_Z8078\: LUT6 
generic map(
  INIT => X"E4E4F0CCCCCCF0CC"
)
port map (
  I0 => cpi_a_cnt(1),
  I1 => rfo1_data1(8),
  I2 => rfo2_data1(8),
  I3 => \GRLFPC20.R.A.RS1\(0),
  I4 => \GRLFPC20.R.A.RS1D\,
  I5 => \GRLFPC20.R.A.ST\,
  O => \GRLFPC20.FPI.OP1\(40));
\GRLFPC20.FPI.OP1[47]_Z8079\: LUT6_L 
generic map(
  INIT => X"E4E4F0CCCCCCF0CC"
)
port map (
  I0 => cpi_a_cnt(1),
  I1 => rfo1_data1(15),
  I2 => rfo2_data1(15),
  I3 => \GRLFPC20.R.A.RS1\(0),
  I4 => \GRLFPC20.R.A.RS1D\,
  I5 => \GRLFPC20.R.A.ST\,
  LO => \GRLFPC20.FPI.OP1\(47));
\GRLFPC20.FPI.OP1[51]_Z8080\: LUT6 
generic map(
  INIT => X"E4E4F0CCCCCCF0CC"
)
port map (
  I0 => cpi_a_cnt(1),
  I1 => rfo1_data1(19),
  I2 => rfo2_data1(19),
  I3 => \GRLFPC20.R.A.RS1\(0),
  I4 => \GRLFPC20.R.A.RS1D\,
  I5 => \GRLFPC20.R.A.ST\,
  O => \GRLFPC20.FPI.OP1\(51));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0[235]_Z8081\: LUT6 
generic map(
  INIT => X"00CC00AAF0F0F0F0"
)
port map (
  I0 => rfo1_data2(29),
  I1 => rfo2_data2(29),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(235),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I4 => \GRLFPC20.COMB.UN1_FPCI_4\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8581\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_RNO[5]\: LUT6 
generic map(
  INIT => X"0000004000000004"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_6095_A2_12_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIOG1B1[91]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(24));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI0UD61[253]\: LUT5 
generic map(
  INIT => X"AAF0CC00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(253),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(240),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIA8LH1[252]\: LUT6 
generic map(
  INIT => X"AAAAF000CCCC0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(252),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(239),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIRM4R[234]\: LUT4 
generic map(
  INIT => X"C0A0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(234),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(247),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(10));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_RNIMQU91[3]\: LUT5 
generic map(
  INIT => X"F0F0EE00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(3),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(5),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(114),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A8_4_0_0[62]\: LUT6 
generic map(
  INIT => X"50000000C0000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1157\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIV0QS[100]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(15));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNITK0B1[87]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(28));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_2_3[13]\: LUT5 
generic map(
  INIT => X"00000020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9551_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_7_TZ[56]_Z8092\: LUT6 
generic map(
  INIT => X"CC44004400000040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_7_TZ\(56));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI5BU51[115]\: LUT5 
generic map(
  INIT => X"AAAAFC00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(115),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(5),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_1[59]_Z8094\: LUT6 
generic map(
  INIT => X"000040400000EA40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9973_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10734\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10767_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_776\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_741\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_1\(59));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A8_5_2[62]_Z8095\: LUT6 
generic map(
  INIT => X"000000000000002B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A8_5_2\(62));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A26_3_1[60]_Z8096\: LUT6_L 
generic map(
  INIT => X"0000A2000000A800"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A26_3_1\(60));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIVN1B1[98]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(17));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIQI1B1[93]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(22));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIPH1B1[92]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(23));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_3_1[32]_Z8100\: LUT6_L 
generic map(
  INIT => X"0000040100000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_3_1\(32));
\GRLFPC20.COMB.V.E.STDATA_1_0[22]\: LUT4 
generic map(
  INIT => X"F2D0"
)
port map (
  I0 => cpi_a_cnt(0),
  I1 => cpi_a_cnt(1),
  I2 => \GRLFPC20.R.I.INST\(22),
  I3 => \GRLFPC20.R.I.PC\(22),
  O => \GRLFPC20.N_2361\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNISJ0B1[86]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(29));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIRI0B1[85]\: LUT4 
generic map(
  INIT => X"ACA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(30));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_9_1[52]_Z8104\: LUT6 
generic map(
  INIT => X"0000000000000080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_9_1\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_6_1[25]_Z8105\: LUT6_L 
generic map(
  INIT => X"0000000000410000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_6_1\(25));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI86LH1[251]\: LUT6 
generic map(
  INIT => X"AAAAF000CCCC0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(251),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(238),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2_RNO[56]\: LUT5 
generic map(
  INIT => X"10000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1012\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_16_TZ[54]_Z8108\: LUT5 
generic map(
  INIT => X"00010088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_16_TZ\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_RNO[61]\: LUT5 
generic map(
  INIT => X"00018000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => N_3105_TZ);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.SIGNRESULT\: LUT5 
generic map(
  INIT => X"0AA019A2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(23),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(24),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(13),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(12),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
  O => \GRLFPC20.FPO.SIGN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_33_RNO\: LUT6 
generic map(
  INIT => X"0F3C2DC30F0F2D0F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(33),
  O => N_3765);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A15_6[18]\: LUT4 
generic map(
  INIT => X"0020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9605\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_5[47]\: LUT6 
generic map(
  INIT => X"A000802000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10088\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_1[52]\: LUT6 
generic map(
  INIT => X"0000000000008020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10225\);
\GRLFPC20.FPI.OP1[36]_Z8115\: LUT6 
generic map(
  INIT => X"E4E4F0CCCCCCF0CC"
)
port map (
  I0 => cpi_a_cnt(1),
  I1 => rfo1_data1(4),
  I2 => rfo2_data1(4),
  I3 => \GRLFPC20.R.A.RS1\(0),
  I4 => \GRLFPC20.R.A.RS1D\,
  I5 => \GRLFPC20.R.A.ST\,
  O => \GRLFPC20.FPI.OP1\(36));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIJTDR1[5]\: LUT6 
generic map(
  INIT => X"0000000200000000"
)
port map (
  I0 => rst,
  I1 => \GRLFPC20.R.MK.LDOP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(5),
  I3 => \GRLFPC20.R.MK.RST\,
  I4 => \GRLFPC20.R.MK.RST2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\);
\GRLFPC20.FPI.OP1[33]_Z8117\: LUT6_L 
generic map(
  INIT => X"E4E4F0CCCCCCF0CC"
)
port map (
  I0 => cpi_a_cnt(1),
  I1 => rfo1_data1(1),
  I2 => rfo2_data1(1),
  I3 => \GRLFPC20.R.A.RS1\(0),
  I4 => \GRLFPC20.R.A.RS1D\,
  I5 => \GRLFPC20.R.A.ST\,
  LO => \GRLFPC20.FPI.OP1\(33));
\GRLFPC20.FPI.OP1[32]_Z8118\: LUT6 
generic map(
  INIT => X"E4E4F0CCCCCCF0CC"
)
port map (
  I0 => cpi_a_cnt(1),
  I1 => rfo1_data1(0),
  I2 => rfo2_data1(0),
  I3 => \GRLFPC20.R.A.RS1\(0),
  I4 => \GRLFPC20.R.A.RS1D\,
  I5 => \GRLFPC20.R.A.ST\,
  O => \GRLFPC20.FPI.OP1\(32));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_0_YY_RNIDKHG3[3]\: LUT6 
generic map(
  INIT => X"55555659A9A6AAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(3),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  I4 => N_6682,
  I5 => N_6683,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_0_YY_RNI47UP3[2]\: LUT6 
generic map(
  INIT => X"55555659A9A6AAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(2),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  I4 => N_6674,
  I5 => N_6675,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_0_YY_RNIBIHG3[4]\: LUT6 
generic map(
  INIT => X"55555659A9A6AAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(4),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  I4 => N_6690,
  I5 => N_6691,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_4\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_Z8122\: LUT6 
generic map(
  INIT => X"0002000200000002"
)
port map (
  I0 => rst,
  I1 => \GRLFPC20.R.MK.LDOP\,
  I2 => \GRLFPC20.R.MK.RST\,
  I3 => \GRLFPC20.R.MK.RST2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14_2\(77),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14\(77),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[37]_Z8123\: LUT6 
generic map(
  INIT => X"FFFFFFFF66F600F0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2630\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_143\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1347\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_972\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0\(37));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15_0_0_O2[39]\: LUT6 
generic map(
  INIT => X"FFFFFFFFFF069000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9389_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1169\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2764\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_782\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1776\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_9[61]\: LUT6 
generic map(
  INIT => X"0000000000080000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_831\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10892\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_9[13]\: LUT6_L 
generic map(
  INIT => X"4800000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9558\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0[18]_Z8127\: LUT6 
generic map(
  INIT => X"FFFFFFFF00200000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10332\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_289\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9604\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(18));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[13]\: LUT5 
generic map(
  INIT => X"FFC43B00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(44),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(48),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8242\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[12]\: LUT5 
generic map(
  INIT => X"FFC43B00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(45),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(49),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8243\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[10]\: LUT5 
generic map(
  INIT => X"FF3BC400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(51),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(47),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8245\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[14]\: LUT5 
generic map(
  INIT => X"FFC43B00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(43),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(47),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8241\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[11]\: LUT5 
generic map(
  INIT => X"FFC43B00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(46),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(50),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8244\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8[9]\: LUT5 
generic map(
  INIT => X"FFC43B00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(48),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(52),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8246\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.NORMDETECT.NOTSLFROMNORM_17_3_0_.M5_I_0\: LUT5 
generic map(
  INIT => X"00010000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_9_REP1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_9\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_93\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M13[1]_Z8135\: LUT5 
generic map(
  INIT => X"55455544"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_3_REP1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M8\(1),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M13\(1));
\GRLFPC20.R.I.INST_RNIHCAM3[19]\: LUT6 
generic map(
  INIT => X"CACCCCCC00000000"
)
port map (
  I0 => cpi_x_inst(19),
  I1 => \GRLFPC20.R.I.INST\(19),
  I2 => \GRLFPC20.R.I.EXEC\,
  I3 => \GRLFPC20.R.I.V\,
  I4 => \GRLFPC20.R.X.FPOP\,
  I5 => \GRLFPC20.N_2146\,
  O => \GRLFPC20.N_1837\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15_0_0[16]_Z8137\: LUT6 
generic map(
  INIT => X"FFFFFFFF28000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2630\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_534\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15_0_0\(16));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_6[6]\: LUT6 
generic map(
  INIT => X"0000020000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9785_1_I_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9497\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1[18]_Z8139\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0001"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10576\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9629\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1034\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_1\(18),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(18));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNO[61]\: LUT6_L 
generic map(
  INIT => X"00000000000000EF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9855_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_3\(60),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_6_2\(60),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2_2\(60),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10788_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A26_20[60]\: LUT6_L 
generic map(
  INIT => X"0000000400000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9508_1\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10839\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0[6]_Z8142\: LUT6_L 
generic map(
  INIT => X"FFFF480048004800"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9664_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9394_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2772\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.TEMP_Z8143\: LUT6 
generic map(
  INIT => X"FFFF0000FFFF2220"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(21),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(77),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(76),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(75),
  I4 => \GRLFPC20.FPI.LDOP\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14\(77),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN_Z8144\: LUT6 
generic map(
  INIT => X"FF000000FF005400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(77),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(76),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(75),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.FPI.LDOP\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14\(77),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.MIFROMINST_Z8145\: LUT6_L 
generic map(
  INIT => X"FFFF0000DDDF0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(63),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(77),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(76),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(75),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.TEMP_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.MIFROMINST\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNISVMB2[63]\: LUT6 
generic map(
  INIT => X"000000002220FFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(63),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(77),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(76),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(75),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.TEMP_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_0_SN_N_6_MUX\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SS0_0\: LUT6 
generic map(
  INIT => X"FFFFFFFFEAC0153F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(9),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(12),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(11),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(374),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SS0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1S2\: LUT6 
generic map(
  INIT => X"FFFFEAC0FFFF153F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(9),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(12),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(11),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(374),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1[6]_Z8149\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF1000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1229\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_291_I\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9511\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9494\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_1[6]_Z8150\: LUT6 
generic map(
  INIT => X"FFFFFFFF003E0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9629\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10025_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1047\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_1\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_8[61]\: LUT6 
generic map(
  INIT => X"0000000000002000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_304\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10891\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_1_LUT6_2_RNI31CV[0]\: LUT5 
generic map(
  INIT => X"AFCFA0C0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(257),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8532\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0[27]_Z8153\: LUT6_L 
generic map(
  INIT => X"FF00FF0006060000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10130\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9509_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9601_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9800_2\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0\(27));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4.Z_AXB1_Z8154\: LUT5 
generic map(
  INIT => X"D22D2DD2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(316),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4.Z_AXB1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_2_RNIKD5I1\: LUT5 
generic map(
  INIT => X"F2002000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(316),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO0_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_2_RNIB1IF5\: LUT6 
generic map(
  INIT => X"FFF2FF20F2002000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(316),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2966_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_RNI5O431\: LUT4 
generic map(
  INIT => X"F220"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(316),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2963_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_61_1.CO0\: LUT6 
generic map(
  INIT => X"0FF2FF2002002000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(316),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_2.CO2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_58_2.ANC1\: LUT6 
generic map(
  INIT => X"0DF2DF2000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(316),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_58_2.CO1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_61_1.SUM0_0_A2\: LUT6 
generic map(
  INIT => X"F20D20DF0DF2DF20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(316),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_61\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"2DD2D22DD22D2DD2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(316),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.SI_63\(50));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2_LUT6_2_RNI7QM32[3]\: LUT6 
generic map(
  INIT => X"FFCEFF0000CE0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8548\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2_LUT6_2_RNIBUM32[7]\: LUT6 
generic map(
  INIT => X"FF08FF0000080000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8552\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_9_RNO\: LUT6 
generic map(
  INIT => X"F0F0F8F000000800"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8554\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(9));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2_LUT6_2_RNICVM32[8]\: LUT6 
generic map(
  INIT => X"FF08FF0000080000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8553\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(8));
\GRLFPC20.COMB.RS1D_1_U\: LUT5_L 
generic map(
  INIT => X"FFBF4000"
)
port map (
  I0 => cpi_d_inst(30),
  I1 => cpi_d_inst(31),
  I2 => \GRLFPC20.N_940\,
  I3 => \GRLFPC20.COMB.FPDECODE.RS1D5\,
  I4 => \GRLFPC20.RS1D_CNST\,
  LO => \GRLFPC20.COMB.RS1D_1\);
\GRLFPC20.UN1_FPOP7_0_A3_0_1\: LUT6 
generic map(
  INIT => X"0000001400000010"
)
port map (
  I0 => cpi_d_inst(9),
  I1 => cpi_d_inst(10),
  I2 => cpi_d_inst(11),
  I3 => cpi_d_inst(12),
  I4 => cpi_d_inst(13),
  I5 => \GRLFPC20.N_3123\,
  O => \GRLFPC20.N_3083_1\);
\GRLFPC20.COMB.RSDECODE.RS1V2_0_A3\: LUT6 
generic map(
  INIT => X"0000000600000000"
)
port map (
  I0 => cpi_d_inst(5),
  I1 => cpi_d_inst(6),
  I2 => cpi_d_inst(9),
  I3 => cpi_d_inst(12),
  I4 => cpi_d_inst(13),
  I5 => \GRLFPC20.N_3117\,
  O => \GRLFPC20.N_3081\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23[113]_Z8169\: LUT6 
generic map(
  INIT => X"5F5F33FF00000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(113));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_Z8170\: LUT6 
generic map(
  INIT => X"53F35FFFFFAFFCAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP[0]_Z8171\: LUT6 
generic map(
  INIT => X"50503300F0F0FF00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_Z8172\: LUT6 
generic map(
  INIT => X"53F35FFFFFAFFCAC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS_LUT6_2_RNIU53L1[4]\: LUT6 
generic map(
  INIT => X"965AF05A3CF05AF0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(234),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(247),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1323\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_10\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS_LUT6_2_RNIS33L1[4]\: LUT6 
generic map(
  INIT => X"965AF05A3CF05AF0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(233),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(246),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1323\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_11\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_1_RNO\: LUT5 
generic map(
  INIT => X"AFCFA0C0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(256),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(243),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8533\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_4_0[56]_Z8176\: LUT6 
generic map(
  INIT => X"DCCC1000CCFF0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10671_I\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1272\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9858_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_4_0\(56));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_2[31]_Z8177\: LUT6 
generic map(
  INIT => X"FFFFFFFF02002200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_76\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10207_I_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_406\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_2_0\(31),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_2\(31));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2[49]_Z8178\: LUT6 
generic map(
  INIT => X"FFFFFFFFDFDD0A00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_715\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2605\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2764\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2161\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2\(49));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_0[42]\: LUT6_L 
generic map(
  INIT => X"0000000000100000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_234\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2220\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15[43]\: LUT6 
generic map(
  INIT => X"0000000000100000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1536_I\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2216\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_0_0_A2[39]\: LUT6 
generic map(
  INIT => X"0000000000000401"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_746\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2233\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_2[36]\: LUT6 
generic map(
  INIT => X"000000B0000000BB"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_406\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10024\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_1[36]_Z8183\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF00001000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9858_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_328\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9971\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_1\(36));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9[27]_Z8184\: LUT6 
generic map(
  INIT => X"4100C3820000C300"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10006\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9972_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9\(27));
\GRLFPC20.COMB.ANNULRES_1_IV_RNO\: LUT6_L 
generic map(
  INIT => X"0000000001000000"
)
port map (
  I0 => cpi_flush,
  I1 => cpi_x_annul,
  I2 => cpi_x_trap,
  I3 => \GRLFPC20.R.X.SEQERR\,
  I4 => \GRLFPC20.N_1494\,
  I5 => \GRLFPC20.N_2015\,
  LO => \GRLFPC20.R.X.SEQERR_M\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[42]_Z8186\: LUT5 
generic map(
  INIT => X"00C43BFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8215\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8213\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(42));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[47]_Z8187\: LUT5 
generic map(
  INIT => X"003BC4FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8208\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8210\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[19]_Z8188\: LUT5 
generic map(
  INIT => X"00C43BFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8238\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8236\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[46]_Z8189\: LUT5 
generic map(
  INIT => X"003BC4FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8209\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8211\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(46));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[50]_Z8190\: LUT5 
generic map(
  INIT => X"003BC4FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8205\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8207\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(50));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[48]_Z8191\: LUT5 
generic map(
  INIT => X"003BC4FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8207\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8209\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(48));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[27]_Z8192\: LUT5 
generic map(
  INIT => X"003BC4FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8228\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8230\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(27));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[39]_Z8193\: LUT5 
generic map(
  INIT => X"00C43BFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8218\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8216\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(39));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[45]_Z8194\: LUT5 
generic map(
  INIT => X"003BC4FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8210\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8212\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(45));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[25]_Z8195\: LUT5 
generic map(
  INIT => X"003BC4FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8230\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8232\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(25));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[52]_Z8196\: LUT5 
generic map(
  INIT => X"00C43BFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8205\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8203\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[53]_Z8197\: LUT5 
generic map(
  INIT => X"00C43BFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8204\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8202\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(53));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[49]_Z8198\: LUT5 
generic map(
  INIT => X"003BC4FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8206\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8208\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(49));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[54]_Z8199\: LUT5 
generic map(
  INIT => X"00C43BFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8203\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8201\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6[51]_Z8200\: LUT5 
generic map(
  INIT => X"00C43BFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8206\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8204\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(51));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[7]_Z8201\: LUT6_L 
generic map(
  INIT => X"000090FF6F00FFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(257),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(7),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(6),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[6]_Z8202\: LUT6_L 
generic map(
  INIT => X"00006F0090FFFFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(257),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(5),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(6),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[4]_Z8203\: LUT6 
generic map(
  INIT => X"00006F0090FFFFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(257),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(4),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[5]_Z8204\: LUT6_L 
generic map(
  INIT => X"00006F0090FFFFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(257),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(4),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(5),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[8]_Z8205\: LUT6_L 
generic map(
  INIT => X"00006F0090FFFFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(257),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(7),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(8),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(8));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10[9]_Z8206\: LUT6_L 
generic map(
  INIT => X"00006F0090FFFFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(257),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(9),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(9));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_12[19]\: LUT6_L 
generic map(
  INIT => X"0040000000400040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_783\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9604_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_717\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9663\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15[28]\: LUT6_L 
generic map(
  INIT => X"0010500000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10860\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2341\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1[41]_Z8209\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFB4000400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_775\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10223_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2707\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2224\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1\(41));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15[42]\: LUT6 
generic map(
  INIT => X"3333333310000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9671_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2842\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2219\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"0DF2DF20F20D20DF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(366),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_457\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.CIN_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.SI_54\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.SI_112\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55.Z_C2_Z8212\: LUT6 
generic map(
  INIT => X"2DFFD2FF002D00D2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(366),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_453\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.CIN_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"D22D2DD22DD2D22D"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(366),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_453\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.CIN_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_113\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48.Z_C2_Z8214\: LUT6 
generic map(
  INIT => X"F2FF20FF00F20020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(360),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(13),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_521\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.SI_48\(9),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"0DF2DF20F20D20DF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(360),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(13),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_521\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.SI_48\(9),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.SI_106\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40.Z_AXBXC0\: LUT4 
generic map(
  INIT => X"2DD2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(352),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(21),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.SI_41\(16));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40.Z_C2_Z8217\: LUT6 
generic map(
  INIT => X"F2FF20FF00F20020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(352),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(21),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_554\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.SI_40\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40.Z_AXBXC1\: LUT6 
generic map(
  INIT => X"0DF2DF20F20D20DF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(352),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(21),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_554\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.CIN_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.SI_40\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.SI_98\(15));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNIEIAI1[28]\: LUT6 
generic map(
  INIT => X"535FACA0ACA0535F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(28),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_28\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNIEIAI1[26]\: LUT6 
generic map(
  INIT => X"535FACA0ACA0535F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(26),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_26\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNIEIAI1[27]\: LUT6 
generic map(
  INIT => X"535FACA0ACA0535F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(27),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_27\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNIEIAI1[29]\: LUT6 
generic map(
  INIT => X"535FACA0ACA0535F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(29),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_29\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNI5ABI1[30]\: LUT6 
generic map(
  INIT => X"535FACA0ACA0535F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(30),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_30\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNICP241[14]\: LUT6 
generic map(
  INIT => X"535FACA0ACA0535F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(14),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_14\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNIEIAI1[19]\: LUT6 
generic map(
  INIT => X"535FACA0ACA0535F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(19),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_19\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNI5ABI1[20]\: LUT6 
generic map(
  INIT => X"535FACA0ACA0535F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(20),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_20\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNI5ABI1[21]\: LUT6 
generic map(
  INIT => X"535FACA0ACA0535F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(21),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_21\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNI5ABI1[25]\: LUT6 
generic map(
  INIT => X"535FACA0ACA0535F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(25),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_25\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNIEIAI1[18]\: LUT6 
generic map(
  INIT => X"535FACA0ACA0535F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(18),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_18\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNI5ABI1[23]\: LUT6 
generic map(
  INIT => X"535FACA0ACA0535F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(23),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_23\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNI5ABI1[24]\: LUT6 
generic map(
  INIT => X"535FACA0ACA0535F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(24),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_24\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNI5ABI1[22]\: LUT6 
generic map(
  INIT => X"535FACA0ACA0535F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(22),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_22\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNICP241[15]\: LUT6 
generic map(
  INIT => X"535FACA0ACA0535F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(15),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_15\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNIEIAI1[17]\: LUT6 
generic map(
  INIT => X"535FACA0ACA0535F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_17\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNIEIAI1[16]\: LUT6 
generic map(
  INIT => X"535FACA0ACA0535F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(16),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_16\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_1_0[47]_Z8236\: LUT6 
generic map(
  INIT => X"5A7B002100000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_796\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9404_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9738_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_1_0\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_O2_0[24]_Z8237\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF00000009"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9785_1_I_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_765\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1231\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_O2_0\(24));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[22]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF1400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9453_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2403\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1775\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(22));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_5_1[60]_Z8239\: LUT6 
generic map(
  INIT => X"00000000C600C644"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9506_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9666_1_I_0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_5_1\(60));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_9[48]\: LUT6 
generic map(
  INIT => X"0000000004000004"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_234\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10164\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20[48]\: LUT6 
generic map(
  INIT => X"00000000F0F0E000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9563_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9508_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10629_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_749\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10154\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_1[49]_Z8242\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFE000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2797\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2645\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(49),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2159\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_1\(49));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[30]_Z8243\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF09000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_406\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9338_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9670_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(30),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0\(30));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A22[53]\: LUT6 
generic map(
  INIT => X"EA5D000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9975_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9670_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10290\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0[20]\: LUT6_L 
generic map(
  INIT => X"F0F0F6F000006600"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2721\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2583\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_742\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1169\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(20));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A24_1[59]\: LUT6 
generic map(
  INIT => X"1000000015000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9576_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9506_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10748\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4[59]_Z8247\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF10000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9503_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9671_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0\(59),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4\(59));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1[42]_Z8248\: LUT6 
generic map(
  INIT => X"FFFFFFFFFF404040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2706\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2724\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10246_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2220\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1\(42));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_11[57]\: LUT6_L 
generic map(
  INIT => X"0000002000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9505_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1230\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10616\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_2[25]\: LUT6 
generic map(
  INIT => X"0250000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9975_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9389_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9719\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2[53]_Z8251\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0004"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12196_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9670_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10305\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10300\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2\(53));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_4[47]_Z8252\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF0020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9492_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_909\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_4_0\(47),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1014\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_4\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_0[11]\: LUT6 
generic map(
  INIT => X"0000000000BA0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10734\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_52\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12250\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_3[11]_Z8254\: LUT6 
generic map(
  INIT => X"FFFFFFFF20000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_751_I\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9858_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_3_0\(11),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_3\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_22[55]\: LUT6 
generic map(
  INIT => X"0010000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9850_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9670_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10460\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_5[6]\: LUT6_L 
generic map(
  INIT => X"0000040000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9700_I\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9496\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0[5]_Z8257\: LUT6 
generic map(
  INIT => X"303000003A300A00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_990_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_6095_A2_12_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_135\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_0[13]\: LUT6_L 
generic map(
  INIT => X"0000000000040002"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_222\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9549\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_4[19]\: LUT6 
generic map(
  INIT => X"0000000000000A22"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9629\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9655\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4[57]_Z8260\: LUT6 
generic map(
  INIT => X"FFFFFFFF00200000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1149\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9670_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10025_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0\(57),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_11[48]\: LUT6 
generic map(
  INIT => X"000000000000A080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_261\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_795\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10166\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0[55]_Z8262\: LUT6_L 
generic map(
  INIT => X"D1FBC0C011BB0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10437_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10624_3\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0\(55));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_9[25]\: LUT6 
generic map(
  INIT => X"0000000000000080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9726\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_3[54]\: LUT6 
generic map(
  INIT => X"0000000000800040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_795\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10365\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_8[55]\: LUT6 
generic map(
  INIT => X"0000000041000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9320_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10410\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10446\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A26_4[56]\: LUT6 
generic map(
  INIT => X"0000000008080008"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9790_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9453_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10524\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2[25]_Z8267\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9748\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_720\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9719\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0\(25),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2\(25));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_0[52]\: LUT6_L 
generic map(
  INIT => X"00D5000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10888_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9394_2\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10224\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4[52]_Z8269\: LUT6 
generic map(
  INIT => X"FFFFFFFF00000008"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9492_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_909\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0\(52),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15[44]\: LUT6_L 
generic map(
  INIT => X"0000000000008020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_909\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_715\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2210\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_1[6]_Z8271\: LUT6 
generic map(
  INIT => X"B888888830000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9665_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9600_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2162_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_1\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_18[33]\: LUT6 
generic map(
  INIT => X"0000000000800000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_328\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9922\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2_0[60]_Z8273\: LUT6 
generic map(
  INIT => X"A0A0B0B000003010"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10767_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12195\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A26_3_1\(60),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2_0\(60));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_19[55]\: LUT6 
generic map(
  INIT => X"0000000004000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9785_1_I_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10457\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_0[36]\: LUT6 
generic map(
  INIT => X"0000000000008C9D"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9828\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_409\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10022\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A26_0[60]\: LUT6 
generic map(
  INIT => X"0000070200000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9671_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10819\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_0_1[60]_Z8277\: LUT6_L 
generic map(
  INIT => X"00FF00000EFF0E0E"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_125\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_746\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10087_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9666_1_I_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_0_1\(60));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_4_0[47]_Z8278\: LUT6 
generic map(
  INIT => X"AB03AA0003030000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10759_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2630\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_4_0\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_20[27]\: LUT6_L 
generic map(
  INIT => X"0000000000000002"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9799\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_4[56]_Z8280\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFE000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1333\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_4_0\(56),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9338\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_4\(56));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0[62]_Z8281\: LUT6_L 
generic map(
  INIT => X"3030743000004400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10917\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1157\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(62));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A22_9[53]\: LUT6_L 
generic map(
  INIT => X"0000000008000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_907\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_304\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10300\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_1[58]_Z8283\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF00200000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_409\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9861_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10678\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_1\(58));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_1[19]_Z8284\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF80F0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9669_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9655\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(19),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_1\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_1[58]_Z8285\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF00080000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10869\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_314_I\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_291_I\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10690\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_1\(58));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_9[19]\: LUT6 
generic map(
  INIT => X"0000000040040000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_796\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9660\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0[19]_Z8287\: LUT6_L 
generic map(
  INIT => X"002000200030A030"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_59\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_796\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNI27BI1[31]\: LUT6 
generic map(
  INIT => X"335FCCA0CCA0335F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(4),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(31),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_31\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_0[57]\: LUT6 
generic map(
  INIT => X"4501000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9969_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10605\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0[0]_Z8290\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF0010"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9435\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9974\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_22[27]\: LUT6 
generic map(
  INIT => X"0000000000000100"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12195\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9801\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A26_11[56]\: LUT6_L 
generic map(
  INIT => X"0000C44000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9492_1\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10531\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0[48]_Z8293\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF00000008"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9560_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9785_1_I_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10155\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0\(48));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1[58]_Z8294\: LUT6_L 
generic map(
  INIT => X"0000000084AC0028"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1019_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_409\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(58));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4[58]_Z8295\: LUT6 
generic map(
  INIT => X"FFFFFFFF08030000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10869\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9861_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_1\(58),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4\(58));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A24_20[59]\: LUT6 
generic map(
  INIT => X"0000000000040000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_776\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10767\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A22_3[53]\: LUT6 
generic map(
  INIT => X"0000000000B00080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_906\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10294\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A22_6[53]\: LUT6_L 
generic map(
  INIT => X"000000000000040C"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_205\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_289\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10297\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_10[55]\: LUT6 
generic map(
  INIT => X"0000000000008808"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9785_1_I_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10448\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A22_8[53]\: LUT6 
generic map(
  INIT => X"0000000000020000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_428\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_907\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10299\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_15[48]\: LUT6 
generic map(
  INIT => X"0080000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10948_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10170\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27[11]\: LUT6 
generic map(
  INIT => X"0000000000C800C0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10734\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9314\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_1[33]_Z8303\: LUT6 
generic map(
  INIT => X"1000100010331000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9896\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9739_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9911_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_328\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_1\(33));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_8[48]\: LUT6_L 
generic map(
  INIT => X"00000000B0100000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9738_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10163\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_4[6]\: LUT6 
generic map(
  INIT => X"0000000100000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9473\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9495\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[54]_Z8306\: LUT6_L 
generic map(
  INIT => X"FF4FB404FB4BB000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(54),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(53),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(52),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[40]_Z8307\: LUT6_L 
generic map(
  INIT => X"FFFBB4B04F4B0400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(38),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(39),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(40),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(40));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[37]_Z8308\: LUT6_L 
generic map(
  INIT => X"FF4FFB4BB404B000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(37),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(35),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(36),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(37));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[52]_Z8309\: LUT6_L 
generic map(
  INIT => X"FFFBB4B04F4B0400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(50),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(51),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(52),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[49]_Z8310\: LUT6_L 
generic map(
  INIT => X"FFB44F04FBB04B00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(48),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(49),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(47),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(49));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[50]_Z8311\: LUT6_L 
generic map(
  INIT => X"FFFBB4B04F4B0400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(48),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(49),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(50),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(50));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[26]_Z8312\: LUT6 
generic map(
  INIT => X"BB0BB000FF4FF444"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(26),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(25),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(25),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(26));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[48]_Z8313\: LUT6_L 
generic map(
  INIT => X"FF4FFB4BB404B000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(48),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(46),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(47),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(48));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[39]_Z8314\: LUT6_L 
generic map(
  INIT => X"FFFBB4B04F4B0400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(37),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(38),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(39),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(39));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[38]_Z8315\: LUT6_L 
generic map(
  INIT => X"FFB44F04FBB04B00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(37),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(38),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(36),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(38));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[47]_Z8316\: LUT6_L 
generic map(
  INIT => X"FFFBB4B04F4B0400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(45),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(46),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(47),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[33]_Z8317\: LUT6_L 
generic map(
  INIT => X"FFFB4F4BB4B00400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(31),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(33),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(32),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(33));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[35]_Z8318\: LUT6_L 
generic map(
  INIT => X"FF4FFB4BB404B000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(35),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(33),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(34),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(35));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[51]_Z8319\: LUT6_L 
generic map(
  INIT => X"FFFBB4B04F4B0400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(49),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(50),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(51),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(51));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[36]_Z8320\: LUT6 
generic map(
  INIT => X"FFB4FBB04F044B00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(35),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(34),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(36),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(36));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[46]_Z8321\: LUT6_L 
generic map(
  INIT => X"BBB00B00FFF44F44"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(45),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(46),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(45),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(46));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[53]_Z8322\: LUT6_L 
generic map(
  INIT => X"FFFB4F4BB4B00400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(51),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(53),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(52),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(53));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[11]_Z8323\: LUT6_L 
generic map(
  INIT => X"FF4FFB4BB404B000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(11),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(9),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(10),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[30]_Z8324\: LUT6 
generic map(
  INIT => X"FFFBB4B04F4B0400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(28),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(29),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(30),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(30));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[10]_Z8325\: LUT6_L 
generic map(
  INIT => X"FFFBB4B04F4B0400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(8),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(9),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(10),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(10));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[42]_Z8326\: LUT6_L 
generic map(
  INIT => X"FF4FFB4BB404B000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(42),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(40),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(41),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(42));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[55]_Z8327\: LUT4_L 
generic map(
  INIT => X"04BF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(54),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(55),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(55));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[34]_Z8328\: LUT6_L 
generic map(
  INIT => X"FFB4FBB04F044B00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(33),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(32),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(34),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(34));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[18]_Z8329\: LUT6 
generic map(
  INIT => X"FFB44F04FBB04B00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(17),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(18),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(16),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(18));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[27]_Z8330\: LUT6 
generic map(
  INIT => X"FFB4FBB04F044B00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(26),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(25),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(27),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(27));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[19]_Z8331\: LUT6 
generic map(
  INIT => X"FF4FFB4BB404B000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(19),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(17),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(18),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[28]_Z8332\: LUT6 
generic map(
  INIT => X"FF4FFB4BB404B000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(28),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(26),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(27),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(28));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[16]_Z8333\: LUT6 
generic map(
  INIT => X"FFFBB4B04F4B0400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(14),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(15),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(16),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(16));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[17]_Z8334\: LUT6 
generic map(
  INIT => X"FF4FFB4BB404B000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(17),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(15),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(16),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(17));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[29]_Z8335\: LUT6 
generic map(
  INIT => X"FFB44F04FBB04B00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(28),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(29),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(27),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(29));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[32]_Z8336\: LUT6_L 
generic map(
  INIT => X"FFB4FBB04F044B00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(31),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(30),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(32),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(32));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[41]_Z8337\: LUT6_L 
generic map(
  INIT => X"FFFBB4B04F4B0400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(39),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(40),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(41),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(41));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[31]_Z8338\: LUT6 
generic map(
  INIT => X"FFFB4F4BB4B00400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(29),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(31),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(30),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(31));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[15]_Z8339\: LUT6_L 
generic map(
  INIT => X"BBB00B00FFF44F44"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_103\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(14),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(15),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(14),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(15));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16[14]_Z8340\: LUT4_L 
generic map(
  INIT => X"0B4F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(14),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(13),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(14));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_4_RNO[47]\: LUT6_L 
generic map(
  INIT => X"0000000001000101"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_715\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_717\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1014\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0[55]_Z8342\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF00000010"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9700_I\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_717\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10456\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(55));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[26]_Z8343\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFFF20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2823\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2379\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2377\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9922\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0\(26));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1[0]_Z8344\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A12_0_0\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9451\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_1\(0),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_5_1[51]_Z8345\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2721\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_0\(51),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2140\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_5_1\(51));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A14_1[34]\: LUT6_L 
generic map(
  INIT => X"0000000000540044"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_751_I\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_720\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12180\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15[12]\: LUT6 
generic map(
  INIT => X"0000000000000102"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_732\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_304\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2475\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_1[50]\: LUT6_L 
generic map(
  INIT => X"0000000000010010"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_909\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2150\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3[55]_Z8349\: LUT6 
generic map(
  INIT => X"FFFFFFFF00CD0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_732\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10479\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0\(55),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3\(55));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15_1_A2[51]\: LUT6 
generic map(
  INIT => X"1010100000100000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2800\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1234\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1650\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[8]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_143\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2584\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2502\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1726\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(8));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_6[7]\: LUT6 
generic map(
  INIT => X"0000000031000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_765\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2512\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15[41]\: LUT6 
generic map(
  INIT => X"0000000012000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2224\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3[6]_Z8354\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9509_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_720\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9495\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0\(6),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_0_RNO[17]\: LUT6 
generic map(
  INIT => X"0000000000080000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9666_1_I_0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_720\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_979\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_0[6]_Z8356\: LUT6 
generic map(
  INIT => X"FFFFFFFFE2000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_0_0\(6),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2563\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_0\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_RNO[5]\: LUT6 
generic map(
  INIT => X"8000808000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1344\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_715\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9861_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_982\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_12[54]_Z8358\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0800"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1169\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8_1\(54),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8_0\(54),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_12\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_4[27]\: LUT6 
generic map(
  INIT => X"44004C0000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10752_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12248\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_8[32]\: LUT6 
generic map(
  INIT => X"0000002800000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9855\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_3[48]\: LUT6 
generic map(
  INIT => X"0000000003000200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9503_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_717\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10158\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_6_0[56]_Z8362\: LUT6_L 
generic map(
  INIT => X"DCCCFCCC10003000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_999_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_795\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1011_1\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_6_0\(56));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_0[51]_Z8363\: LUT6 
generic map(
  INIT => X"F0F0F4F000004400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10746_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2669\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_289\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2594\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_0\(51));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_0[4]_Z8364\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF20000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2645\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9495\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_0\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A22_18[53]\: LUT6 
generic map(
  INIT => X"0000000000000100"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9785_1_I_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10309\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_RNO[13]\: LUT6 
generic map(
  INIT => X"000000000020008A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_202\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9666_1_I_0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1133\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1[62]_Z8367\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A8_5_2\(62),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10926\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10929\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(62),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(62));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2[4]_Z8368\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2772\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2400\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9726\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_0\(4),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_0[36]_Z8369\: LUT6 
generic map(
  INIT => X"FF000000FF001000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12021_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10030_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_328\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_0\(36));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_0[54]_Z8370\: LUT6_L 
generic map(
  INIT => X"D951880051510000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9321_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10383_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9394_2\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_0\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A12_7[0]\: LUT6 
generic map(
  INIT => X"0000000000000010"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9453\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_RNO[5]\: LUT6_L 
generic map(
  INIT => X"0000000010000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_776\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9666_1_I_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_983\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_15[27]\: LUT6 
generic map(
  INIT => X"0000040000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9794\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_13[52]\: LUT6_L 
generic map(
  INIT => X"0000000000100040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_749\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10237\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_2[17]\: LUT6 
generic map(
  INIT => X"0000000020000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9700_I\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2445\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_1[56]_Z8376\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF00001050"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_795\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_328\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_1_0\(56),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_1\(56));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_0[32]_Z8377\: LUT6 
generic map(
  INIT => X"8080001000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9790_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9610_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_0\(32));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A15_5[18]\: LUT6 
generic map(
  INIT => X"0000000088008000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_732\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9604\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0[59]_Z8379\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF00020000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10824_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10456\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(59));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_10[19]\: LUT6 
generic map(
  INIT => X"00000000008C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_775\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9661\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_1_0[31]_Z8381\: LUT6_L 
generic map(
  INIT => X"FA000000FE330000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9797_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10207_I_2\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_796\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_1_0\(31));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15[26]\: LUT6 
generic map(
  INIT => X"0000000000000006"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_717\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2377\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_1[49]_Z8383\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF00000002"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_742\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2167\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_1\(49));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2[28]_Z8384\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0010"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2697\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(28),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(28),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2\(28));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15[43]\: LUT6 
generic map(
  INIT => X"FFFFFFFF00000002"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2214\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1653\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7_1[52]_Z8386\: LUT6 
generic map(
  INIT => X"FFFFFFFF10110000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10207_I_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_909\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10223_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2129\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7_1\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIPN2P1[79]\: LUT5 
generic map(
  INIT => X"00000001"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1006_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_5_RNO[56]\: LUT6 
generic map(
  INIT => X"0000000000040005"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1009\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A15_11_2_I_O2_LUT6_2_RNI4G0G2[18]\: LUT6 
generic map(
  INIT => X"0000000000000001"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2403\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_1[26]\: LUT6 
generic map(
  INIT => X"0000000400000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10948_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9861_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2379\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0[58]_Z8391\: LUT6_L 
generic map(
  INIT => X"0A0A0A0B00000001"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_76\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1019_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A30_10_1\(58),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(58));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_1[5]_Z8392\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF05040000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2608\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1725\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_1\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1[23]_Z8393\: LUT6 
generic map(
  INIT => X"0000000010101110"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(23));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0[28]_Z8394\: LUT6 
generic map(
  INIT => X"0303070300000500"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10891_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2707\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(28));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_0[27]\: LUT6 
generic map(
  INIT => X"00000000400040C0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_289\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9779\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_0_0[31]_Z8396\: LUT6_L 
generic map(
  INIT => X"00008080005580D5"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1553_I\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10790\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_409\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9666_1_I_0\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_0_0\(31));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_4[57]\: LUT6 
generic map(
  INIT => X"C800080000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10943\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10609\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0[33]_Z8398\: LUT6_L 
generic map(
  INIT => X"000000F0008800F8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_23_0\(47),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_328\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_720\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(33));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A15_11_2_I_O2_LUT6_2_RNIDC5P1[18]\: LUT6 
generic map(
  INIT => X"0000000000200000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_989\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15[9]\: LUT6 
generic map(
  INIT => X"0000000040000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2502\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_11[55]\: LUT6 
generic map(
  INIT => X"004C000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1344\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10449\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0[19]_Z8402\: LUT6_L 
generic map(
  INIT => X"0000000072225000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9739_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9642\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9671_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_717\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0[25]_Z8403\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF02C40000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_6095_A2_11_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9726\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0\(25));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_1[28]_Z8404\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF0200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_289\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10246_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2343\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1593\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_1\(28));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27[47]\: LUT6 
generic map(
  INIT => X"0000020002000200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_796\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10082\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0[6]_Z8406\: LUT6 
generic map(
  INIT => X"FFFFFFFF02000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9496\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_9[24]\: LUT6_L 
generic map(
  INIT => X"0000200000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10948_1\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1231\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_4_A2_0_A2[17]\: LUT6 
generic map(
  INIT => X"0000000000000200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_289\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2447\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_5_0_A2[17]\: LUT6 
generic map(
  INIT => X"0002000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10948_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9861_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2448\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIGD5I3[80]\: LUT6 
generic map(
  INIT => X"0000000000020000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10948_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1041\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_3_0[11]_Z8411\: LUT6_L 
generic map(
  INIT => X"CC00800000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9321_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9858_1\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_3_0\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A26_2[56]\: LUT6_L 
generic map(
  INIT => X"5100110000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9858_1\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10522\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_13[11]_Z8413\: LUT6_L 
generic map(
  INIT => X"0000CC0000000400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_125\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1019_1\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_13\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7[55]_Z8414\: LUT6 
generic map(
  INIT => X"FFFFFFFF01020000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1175\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10699\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7\(55));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_6[27]\: LUT6 
generic map(
  INIT => X"0000000020001000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_783\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_909\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9785\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0[15]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFF80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10243_3\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_989\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0\(15),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1725\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(15));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_1[23]\: LUT5 
generic map(
  INIT => X"00800000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1336\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2400\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0[52]_Z8418\: LUT6_L 
generic map(
  INIT => X"B3A0A0A033000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_16_0\(52),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10243_3\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_RNO_0[17]\: LUT6_L 
generic map(
  INIT => X"0000000000000104"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_978\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_2[49]\: LUT6_L 
generic map(
  INIT => X"0000000000080040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12132\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2161\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_0[35]\: LUT6 
generic map(
  INIT => X"000000D000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2584\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2255\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_O2[29]\: LUT6 
generic map(
  INIT => X"0A0A4E0A00004400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1267\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_135\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1342\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_866\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_3[27]\: LUT6_L 
generic map(
  INIT => X"0000000000004004"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9782\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_7[27]\: LUT6_L 
generic map(
  INIT => X"0000000000008880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9786\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_M_RNO[6]\: LUT6 
generic map(
  INIT => X"FFFFDFFF0000D0FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14\(77),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN3_NOTRESETORUNIMP\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8115\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_11\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1[44]_Z8426\: LUT6 
generic map(
  INIT => X"00FF20FF00002020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1011_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12131\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1342\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(44));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_1[55]_Z8427\: LUT6 
generic map(
  INIT => X"0000109000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9850_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_314_I\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_1\(55));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_3[25]\: LUT6 
generic map(
  INIT => X"0000000000200000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10146\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9748\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9720\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A22_1[53]\: LUT6 
generic map(
  INIT => X"7A00000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1149\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_314_I\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10292\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A30_0[58]\: LUT6 
generic map(
  INIT => X"0041000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9861_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10678\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_0[31]_Z8431\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF0000005C"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10006\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_234\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_0_0\(31),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_0\(31));
\GRLFPC20.COMB.V.E.STDATA_1[5]_Z8432\: LUT6_L 
generic map(
  INIT => X"F2D0FFFFF2D00000"
)
port map (
  I0 => cpi_a_cnt(0),
  I1 => cpi_a_cnt(1),
  I2 => \GRLFPC20.R.I.INST\(5),
  I3 => \GRLFPC20.R.I.PC\(5),
  I4 => \GRLFPC20.R.A.AFQ\,
  I5 => \GRLFPC20.N_2377\,
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(5));
\GRLFPC20.COMB.V.E.STDATA_1[3]_Z8433\: LUT6_L 
generic map(
  INIT => X"F2D0FFFFF2D00000"
)
port map (
  I0 => cpi_a_cnt(0),
  I1 => cpi_a_cnt(1),
  I2 => \GRLFPC20.R.I.INST\(3),
  I3 => \GRLFPC20.R.I.PC\(3),
  I4 => \GRLFPC20.R.A.AFQ\,
  I5 => \GRLFPC20.N_2375\,
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(3));
\GRLFPC20.COMB.V.E.STDATA_1[31]_Z8434\: LUT6_L 
generic map(
  INIT => X"F2D0FFFFF2D00000"
)
port map (
  I0 => cpi_a_cnt(0),
  I1 => cpi_a_cnt(1),
  I2 => \GRLFPC20.R.I.INST\(31),
  I3 => \GRLFPC20.R.I.PC\(31),
  I4 => \GRLFPC20.R.A.AFQ\,
  I5 => \GRLFPC20.N_2403\,
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(31));
\GRLFPC20.COMB.V.E.STDATA_1[10]_Z8435\: LUT6_L 
generic map(
  INIT => X"F2D0FFFFF2D00000"
)
port map (
  I0 => cpi_a_cnt(0),
  I1 => cpi_a_cnt(1),
  I2 => \GRLFPC20.R.I.INST\(10),
  I3 => \GRLFPC20.R.I.PC\(10),
  I4 => \GRLFPC20.R.A.AFQ\,
  I5 => \GRLFPC20.N_2382\,
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(10));
\GRLFPC20.COMB.V.E.STDATA_1[2]_Z8436\: LUT6_L 
generic map(
  INIT => X"F2D0FFFFF2D00000"
)
port map (
  I0 => cpi_a_cnt(0),
  I1 => cpi_a_cnt(1),
  I2 => \GRLFPC20.R.I.INST\(2),
  I3 => \GRLFPC20.R.I.PC\(2),
  I4 => \GRLFPC20.R.A.AFQ\,
  I5 => \GRLFPC20.N_2374\,
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(2));
\GRLFPC20.COMB.V.E.STDATA_1[14]_Z8437\: LUT6_L 
generic map(
  INIT => X"F2D0FFFFF2D00000"
)
port map (
  I0 => cpi_a_cnt(0),
  I1 => cpi_a_cnt(1),
  I2 => \GRLFPC20.R.I.INST\(14),
  I3 => \GRLFPC20.R.I.PC\(14),
  I4 => \GRLFPC20.R.A.AFQ\,
  I5 => \GRLFPC20.N_2386\,
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(14));
\GRLFPC20.COMB.V.E.STDATA_1[7]_Z8438\: LUT6_L 
generic map(
  INIT => X"F2D0FFFFF2D00000"
)
port map (
  I0 => cpi_a_cnt(0),
  I1 => cpi_a_cnt(1),
  I2 => \GRLFPC20.R.I.INST\(7),
  I3 => \GRLFPC20.R.I.PC\(7),
  I4 => \GRLFPC20.R.A.AFQ\,
  I5 => \GRLFPC20.N_2379\,
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(7));
\GRLFPC20.COMB.V.E.STDATA_1[13]_Z8439\: LUT6_L 
generic map(
  INIT => X"F2D0FFFFF2D00000"
)
port map (
  I0 => cpi_a_cnt(0),
  I1 => cpi_a_cnt(1),
  I2 => \GRLFPC20.R.I.INST\(13),
  I3 => \GRLFPC20.R.I.PC\(13),
  I4 => \GRLFPC20.R.A.AFQ\,
  I5 => \GRLFPC20.N_2385\,
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(13));
\GRLFPC20.COMB.V.E.STDATA_1[16]_Z8440\: LUT6_L 
generic map(
  INIT => X"F2D0FFFFF2D00000"
)
port map (
  I0 => cpi_a_cnt(0),
  I1 => cpi_a_cnt(1),
  I2 => \GRLFPC20.R.I.INST\(16),
  I3 => \GRLFPC20.R.I.PC\(16),
  I4 => \GRLFPC20.R.A.AFQ\,
  I5 => \GRLFPC20.N_2388\,
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(16));
\GRLFPC20.COMB.V.E.STDATA_1[25]_Z8441\: LUT6_L 
generic map(
  INIT => X"FD20FFFFFD200000"
)
port map (
  I0 => cpi_a_cnt(0),
  I1 => cpi_a_cnt(1),
  I2 => \GRLFPC20.R.I.PC\(25),
  I3 => \GRLFPC20.R.I.INST\(25),
  I4 => \GRLFPC20.R.A.AFQ\,
  I5 => \GRLFPC20.N_2397\,
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(25));
\GRLFPC20.COMB.V.E.STDATA_1[23]_Z8442\: LUT6_L 
generic map(
  INIT => X"F2D0FFFFF2D00000"
)
port map (
  I0 => cpi_a_cnt(0),
  I1 => cpi_a_cnt(1),
  I2 => \GRLFPC20.R.I.INST\(23),
  I3 => \GRLFPC20.R.I.PC\(23),
  I4 => \GRLFPC20.R.A.AFQ\,
  I5 => \GRLFPC20.N_2395\,
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(23));
\GRLFPC20.COMB.V.E.STDATA_1[24]_Z8443\: LUT6_L 
generic map(
  INIT => X"F2D0FFFFF2D00000"
)
port map (
  I0 => cpi_a_cnt(0),
  I1 => cpi_a_cnt(1),
  I2 => \GRLFPC20.R.I.INST\(24),
  I3 => \GRLFPC20.R.I.PC\(24),
  I4 => \GRLFPC20.R.A.AFQ\,
  I5 => \GRLFPC20.N_2396\,
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(24));
\GRLFPC20.COMB.V.E.STDATA_1[27]_Z8444\: LUT6_L 
generic map(
  INIT => X"FD20FFFFFD200000"
)
port map (
  I0 => cpi_a_cnt(0),
  I1 => cpi_a_cnt(1),
  I2 => \GRLFPC20.R.I.PC\(27),
  I3 => \GRLFPC20.R.I.INST\(27),
  I4 => \GRLFPC20.R.A.AFQ\,
  I5 => \GRLFPC20.N_2399\,
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(27));
\GRLFPC20.COMB.V.E.STDATA_1[26]_Z8445\: LUT6_L 
generic map(
  INIT => X"FD20FFFFFD200000"
)
port map (
  I0 => cpi_a_cnt(0),
  I1 => cpi_a_cnt(1),
  I2 => \GRLFPC20.R.I.PC\(26),
  I3 => \GRLFPC20.R.I.INST\(26),
  I4 => \GRLFPC20.R.A.AFQ\,
  I5 => \GRLFPC20.N_2398\,
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(26));
\GRLFPC20.COMB.V.E.STDATA_1[11]_Z8446\: LUT6_L 
generic map(
  INIT => X"F2D0FFFFF2D00000"
)
port map (
  I0 => cpi_a_cnt(0),
  I1 => cpi_a_cnt(1),
  I2 => \GRLFPC20.R.I.INST\(11),
  I3 => \GRLFPC20.R.I.PC\(11),
  I4 => \GRLFPC20.R.A.AFQ\,
  I5 => \GRLFPC20.N_2383\,
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(11));
\GRLFPC20.COMB.V.E.STDATA_1[9]_Z8447\: LUT6_L 
generic map(
  INIT => X"F2D0FFFFF2D00000"
)
port map (
  I0 => cpi_a_cnt(0),
  I1 => cpi_a_cnt(1),
  I2 => \GRLFPC20.R.I.INST\(9),
  I3 => \GRLFPC20.R.I.PC\(9),
  I4 => \GRLFPC20.R.A.AFQ\,
  I5 => \GRLFPC20.N_2381\,
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(9));
\GRLFPC20.COMB.V.E.STDATA_1[4]_Z8448\: LUT6_L 
generic map(
  INIT => X"F2D0FFFFF2D00000"
)
port map (
  I0 => cpi_a_cnt(0),
  I1 => cpi_a_cnt(1),
  I2 => \GRLFPC20.R.I.INST\(4),
  I3 => \GRLFPC20.R.I.PC\(4),
  I4 => \GRLFPC20.R.A.AFQ\,
  I5 => \GRLFPC20.N_2376\,
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(4));
\GRLFPC20.COMB.V.E.STDATA_1[30]_Z8449\: LUT6_L 
generic map(
  INIT => X"F2D0FFFFF2D00000"
)
port map (
  I0 => cpi_a_cnt(0),
  I1 => cpi_a_cnt(1),
  I2 => \GRLFPC20.R.I.INST\(30),
  I3 => \GRLFPC20.R.I.PC\(30),
  I4 => \GRLFPC20.R.A.AFQ\,
  I5 => \GRLFPC20.N_2402\,
  LO => \GRLFPC20.COMB.V.E.STDATA_1\(30));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20[32]\: LUT6 
generic map(
  INIT => X"0000000000066600"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10661\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9846\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_12[48]\: LUT6 
generic map(
  INIT => X"0000000000000084"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_717\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10167\);
\GRLFPC20.COMB.UN4_LOCK\: LUT6 
generic map(
  INIT => X"FFFFFFFFFEFFFEFE"
)
port map (
  I0 => cpi_d_annul,
  I1 => cpi_d_trap,
  I2 => cpi_flush,
  I3 => \GRLFPC20.R.STATE\(1),
  I4 => \GRLFPC20.R.STATE\(0),
  I5 => \GRLFPC20.COMB.LOCKGEN.LOCKI\,
  O => \GRLFPC20.N_1317\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0[32]_Z8453\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0800"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9863_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_0\(32),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9855\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0\(32));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15[28]\: LUT6 
generic map(
  INIT => X"FFFFFFFF08000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2601\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2206\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1593\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_5_A2_0_A2[56]\: LUT6 
generic map(
  INIT => X"0000000000800000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2764\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN[0]_Z8456\: LUT6 
generic map(
  INIT => X"F1F7F1F700F5F5FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(371),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(373),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN3_GEN_0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN1_NOTPROP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8_0_0[57]_Z8457\: LUT6 
generic map(
  INIT => X"FBFBF7F70EFDFD0E"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(371),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(373),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(2),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN1_NOTPROP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8_0_0\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0[13]_Z8458\: LUT6 
generic map(
  INIT => X"8000030380000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_9_0\(25),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A26_22_0\(60),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(13));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_1[29]\: LUT6 
generic map(
  INIT => X"4000000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9861_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2337\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0[3]_Z8460\: LUT6 
generic map(
  INIT => X"FFFFFFFFD8000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10860\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1006\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_1[19]\: LUT6 
generic map(
  INIT => X"0027000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9652_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9652\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13[61]\: LUT6_L 
generic map(
  INIT => X"0000000004030000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10767_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10882\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2_LUT6_2_RNI5T892[3]\: LUT6 
generic map(
  INIT => X"C9C33933363CC6CC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8549\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(4),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_AXB_4\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_3[11]\: LUT6_L 
generic map(
  INIT => X"0000004700000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9858_1\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9318\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_7[47]\: LUT6 
generic map(
  INIT => X"0000000000800000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9296_I\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10090\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_8[51]\: LUT6 
generic map(
  INIT => X"0001000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10943\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2140\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A14_9[34]\: LUT6 
generic map(
  INIT => X"0200000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9974\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_8[11]\: LUT6 
generic map(
  INIT => X"000000008800A000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_742\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9323\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_1[11]\: LUT6 
generic map(
  INIT => X"0222002200000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9330_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9316\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_5[57]\: LUT6 
generic map(
  INIT => X"0000050400000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10943\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12238\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0[34]_Z8471\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0800"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9993\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9974\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(34),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(34));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_11[11]\: LUT6_L 
generic map(
  INIT => X"0100020000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9858_1\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9326\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_38_0[0]\: LUT6_L 
generic map(
  INIT => X"AAAAAAAAAAAACAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(13),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(12),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9249\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_1[48]\: LUT6_L 
generic map(
  INIT => X"000000000004000A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_135\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10156\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A15_11_2_I_O2_LUT6_2_RNIFE5P1[18]\: LUT6 
generic map(
  INIT => X"0000000000000004"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_967\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_10_A2_0_A2[61]\: LUT6 
generic map(
  INIT => X"0000000100000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2762\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_8[49]\: LUT6 
generic map(
  INIT => X"0000000000040000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2167\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_0[20]\: LUT6 
generic map(
  INIT => X"0000004000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9861_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2125\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_5_0[51]_Z8479\: LUT6 
generic map(
  INIT => X"0000440A00000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10157_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_5_0\(51));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_0_1_LUT6_2_RNI156P1[6]\: LUT6 
generic map(
  INIT => X"4000000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9861_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1025\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15[8]\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF4C00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1006_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2448\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_989\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1726\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIAEF42[78]\: LUT6 
generic map(
  INIT => X"0000000000000004"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_991_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_0_1_LUT6_2_RNIU16P1[6]\: LUT6 
generic map(
  INIT => X"0000120000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9861_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1039\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15_1[17]\: LUT6 
generic map(
  INIT => X"FFFFFFFF00000020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_595\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2208\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1710\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5[13]_Z8485\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFFFF40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_8_1\(13),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12249\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1133\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2\(13),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5\(13));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1[29]\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF4440"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1169\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_789\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(29),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_0\(29),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRLOI\(29));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_1[0]_Z8487\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF10000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9916_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9454\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_1\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2[4]\: LUT6 
generic map(
  INIT => X"1000000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2831\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_1[46]\: LUT6 
generic map(
  INIT => X"0000000001000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_921\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2208\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A12_5[0]\: LUT6 
generic map(
  INIT => X"0000000001000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9451\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2[12]\: LUT6 
generic map(
  INIT => X"0000000002000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2842\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_6[57]\: LUT6 
generic map(
  INIT => X"0010000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2730\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A30_21[58]\: LUT6 
generic map(
  INIT => X"0010000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10699\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_57_Z8494\: LUT5 
generic map(
  INIT => X"41B1BE4E"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(57),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_57\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNIU1N42[42]\: LUT6 
generic map(
  INIT => X"65A9CF039A5630FC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(42),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_42\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNIU1N42[52]\: LUT6 
generic map(
  INIT => X"65A9CF039A5630FC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(52),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_52\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNIU1N42[43]\: LUT6 
generic map(
  INIT => X"65A9CF039A5630FC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(43),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_43\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNIU1N42[53]\: LUT6 
generic map(
  INIT => X"65A9CF039A5630FC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(53),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_53\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNIU1N42[51]\: LUT6 
generic map(
  INIT => X"65A9CF039A5630FC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(51),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_51\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNI7AM42[48]\: LUT6 
generic map(
  INIT => X"65A9CF039A5630FC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(48),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_48\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNIU1N42[50]\: LUT6 
generic map(
  INIT => X"65A9CF039A5630FC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(50),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_50\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNI7AM42[49]\: LUT6 
generic map(
  INIT => X"65A9CF039A5630FC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(49),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_49\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNI7AM42[47]\: LUT6 
generic map(
  INIT => X"65A9CF039A5630FC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(47),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_47\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNI7AM42[46]\: LUT6 
generic map(
  INIT => X"65A9CF039A5630FC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(46),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_46\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNIU1N42[45]\: LUT6 
generic map(
  INIT => X"65A9CF039A5630FC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(45),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_45\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNIU1N42[44]\: LUT6 
generic map(
  INIT => X"65A9CF039A5630FC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(44),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_44\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNIU1N42[41]\: LUT6 
generic map(
  INIT => X"65A9CF039A5630FC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(41),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_41\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNIU1N42[40]\: LUT6 
generic map(
  INIT => X"65A9CF039A5630FC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(40),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_40\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNI7AM42[39]\: LUT6 
generic map(
  INIT => X"65A9CF039A5630FC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(39),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_39\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_RNIU1N42[32]\: LUT6 
generic map(
  INIT => X"65A9CF039A5630FC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(32),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_32\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_36_RNO\: LUT6 
generic map(
  INIT => X"0F3C2DC30F0F2D0F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(36),
  O => N_3768);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_54_RNO\: LUT6 
generic map(
  INIT => X"0F3C2DC30F0F2D0F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(54),
  O => N_3786);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_37_RNO\: LUT6 
generic map(
  INIT => X"0F3C2DC30F0F2D0F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(37),
  O => N_3769);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_35_RNO\: LUT6 
generic map(
  INIT => X"0F3C2DC30F0F2D0F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(35),
  O => N_3767);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_38_RNO\: LUT6 
generic map(
  INIT => X"0F3C2DC30F0F2D0F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(38),
  O => N_3770);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_34_RNO\: LUT6 
generic map(
  INIT => X"0F3C2DC30F0F2D0F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(34),
  O => N_3766);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CRY_56_RNO\: LUT6 
generic map(
  INIT => X"0F3C2DC30F0F2D0F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M0\(56),
  O => N_3788);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI8CF42[78]\: LUT6 
generic map(
  INIT => X"0000000000000002"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1006\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O2_3_O2[29]\: LUT6 
generic map(
  INIT => X"0200400012124000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_789\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15[44]\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF8000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2708\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2734\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2140\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1748\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_2[48]\: LUT6 
generic map(
  INIT => X"2100200000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10157_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10157\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3[50]_Z8522\: LUT6 
generic map(
  INIT => X"4A4040400A000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9506_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2600\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2505_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3\(50));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_4_1[31]_Z8523\: LUT6 
generic map(
  INIT => X"00000000010001FA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_406\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10410\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_4_1\(31));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0[53]_Z8524\: LUT6 
generic map(
  INIT => X"0808190800001100"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A22_16_0\(53),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_304\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A22_2_0\(53),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0_0\(53));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1[24]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF1000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9453_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1_0\(24),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1775\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(24));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0[14]_Z8526\: LUT6_L 
generic map(
  INIT => X"FFFFFFFF04000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2454_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2129\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0\(14));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7[48]_Z8527\: LUT6 
generic map(
  INIT => X"FFFFFFFFFFFF1000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_5_0\(48),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2166\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_0\(48),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7\(48));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_0[27]_Z8528\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFD9004000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2517_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9788_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(27),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_0\(27));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2_0[47]_Z8529\: LUT6 
generic map(
  INIT => X"0222002000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9790_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9652_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2_0\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A8_0[62]\: LUT6 
generic map(
  INIT => X"1088000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9655_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9492_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10926\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0[58]_Z8531\: LUT6 
generic map(
  INIT => X"0A001E140A000A00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A30_14_0\(58),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_409\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9558_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_2_0\(58));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A14[34]\: LUT6 
generic map(
  INIT => X"0000406100000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12132\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9738_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9964\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0[49]_Z8533\: LUT6 
generic map(
  INIT => X"5500550000004000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_222\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1283\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_0\(49));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_7[60]_Z8534\: LUT6 
generic map(
  INIT => X"4060406040600000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9652_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10860\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_7\(60));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0[27]_Z8535\: LUT6_L 
generic map(
  INIT => X"02B2000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9601_2\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3_0\(27));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_5_0[11]_Z8536\: LUT6 
generic map(
  INIT => X"0040000000003000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9604_1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_5_0\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A12[0]\: LUT6 
generic map(
  INIT => X"3304300100000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A12_0\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9445\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIM5RH2[226]\: LUT6 
generic map(
  INIT => X"FF000FF033CC55AA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(226),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_5_N_4_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SS0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_5\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST_RNIK6F21[17]\: LUT5 
generic map(
  INIT => X"E2C01D3F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_5_N_4_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIR9QH2[225]\: LUT6 
generic map(
  INIT => X"FF0033CC0FF055AA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(225),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_6_N_4_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SS0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_6\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST_RNISDE21[17]\: LUT5 
generic map(
  INIT => X"E2C01D3F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_6_N_4_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI0EPH2[224]\: LUT6 
generic map(
  INIT => X"FF000FF033CC55AA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(224),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_7_N_4_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SS0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_7\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST_RNIRCE21[17]\: LUT5 
generic map(
  INIT => X"E2C01D3F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_7_N_4_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI6IOH2[223]\: LUT6 
generic map(
  INIT => X"FF0033CC0FF055AA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(223),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_8_N_4_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SS0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_8\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST_RNIRBE21[17]\: LUT5 
generic map(
  INIT => X"D8882777"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(17),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_8_N_4_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIJUOL2[222]\: LUT6 
generic map(
  INIT => X"FF0033CC0FF055AA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(222),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_9_N_4_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SS0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_9\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIBRE61[106]\: LUT5 
generic map(
  INIT => X"ACA0535F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_9_N_4_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIFQOL2[221]\: LUT6 
generic map(
  INIT => X"FF000FF033CC55AA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(221),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_10_N_4_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SS0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_10\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIAQE61[105]\: LUT5 
generic map(
  INIT => X"ACA0535F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_10_N_4_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIBMOL2[220]\: LUT6 
generic map(
  INIT => X"FF0033CC0FF055AA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(220),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_11_N_4_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SS0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_11\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI9PE61[104]\: LUT5 
generic map(
  INIT => X"ACA0535F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_11_N_4_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIGQNL2[219]\: LUT6 
generic map(
  INIT => X"FF000FF033CC55AA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(219),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_12_N_4_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SS0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_12\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI8OE61[103]\: LUT5 
generic map(
  INIT => X"ACA0535F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_12_N_4_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNICMNL2[218]\: LUT6 
generic map(
  INIT => X"FF0033CC0FF055AA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(218),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_13_N_4_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SS0\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SM0\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_13\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI7NE61[102]\: LUT5 
generic map(
  INIT => X"ACA0535F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_13_N_4_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_39_U[0]\: LUT6 
generic map(
  INIT => X"CCCCCCCCAAF0CCF0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(13),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(12),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9257\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_39_U_N_3_3\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_39_U_N_4_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(67),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9260\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_39_U_N_4L6\: LUT4 
generic map(
  INIT => X"00EC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(27),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_39_U_N_4_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M12_RNI0OR65[1]\: LUT6 
generic map(
  INIT => X"E0E0FFE0FCECFFFC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M13\(1),
  I2 => N_14234,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M12\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_I_I_A2_0_O2_1\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_SM12\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.EXPYBUS_1_I_A2_I_RNI0A1V1[1]\: LUT6 
generic map(
  INIT => X"FA00FA300A000A30"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(243),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_584\,
  O => N_14234);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15_FAST[16]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFF1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_135\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_765\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2233\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2156\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15_0_0\(16),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15_1\(16),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_FAST\(16));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST[10]\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(16),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_FAST\(16),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15_REP1[16]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFF1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_135\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_765\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2233\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2156\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15_0_0\(16),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15_1\(16),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_REP1\(16));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_10_REP1\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP1\,
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_REP1\(16),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15_REP2[16]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFF1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_135\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_765\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2233\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2156\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15_0_0\(16),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15_1\(16),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_REP2\(16));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_10_REP2\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_16_REP2\,
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_REP2\(16),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST_RNO[11]\: LUT3_L 
generic map(
  INIT => X"01"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2502\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_2_1\(11),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_7\(11),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9288_I_FAST\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST[11]_Z8570\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(11),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9288_I_FAST\,
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST[9]_Z8571\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(9),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_FAST\(9),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_FAST[374]_Z8572\: LUT5_L 
generic map(
  INIT => X"01FFFF40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_2\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(0),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_FAST\(374));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_FAST[12]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFA8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10157_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2774\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1283\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2337\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1661\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3\(12),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_FAST\(12));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST[12]_Z8574\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(12),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_FAST\(12),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_FAST[1]\: LUT6_L 
generic map(
  INIT => X"FFF2F0F20F020002"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(117),
  I1 => \GRLFPC20.FPI.LDOP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7740\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7976\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_FAST\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_DIVMULTV_FAST[0]_Z8576\: LUT4_L 
generic map(
  INIT => X"4002"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(3),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(2),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF\(0),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_DIVMULTV_FAST\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_FAST[3]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7914\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7738\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7974\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_FAST\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_REP1[3]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7914\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7738\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7974\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_REP1\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_FAST[15]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7902\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7726\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7962\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_FAST\(15));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_FAST[17]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7900\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7724\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7960\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_FAST\(17));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_FAST[8]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7909\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7733\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7969\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_FAST\(8));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_REP1[8]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7909\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7733\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7969\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_REP1\(8));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_FAST[8]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFF0400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_143\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2584\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2502\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1726\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_FAST\(8));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST[8]_Z8584\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(8),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_FAST\(8),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_FAST[19]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_0\(19),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_5_1\(19),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4\(19),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8\(19),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7\(19),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6\(19),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_FAST\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST[19]_Z8586\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(19),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_FAST\(19),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST[29]_Z8587\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(29),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRLOI\(29),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_29_REP1_Z8588\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_29_REP1\,
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRLOI\(29),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST[30]_Z8589\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(30),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRLOI\(30),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_30_REP1_Z8590\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_30_REP1\,
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRLOI\(30),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_FAST[17]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1711\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1648\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1710\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_0\(17),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1661\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_1\(17),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_FAST\(17));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST[17]_Z8592\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(17),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_FAST\(17),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_REP1[17]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1711\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1648\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1710\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_0\(17),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1661\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_1\(17),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_REP1\(17));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP1_Z8594\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP1\,
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_REP1\(17),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_REP2[17]\: LUT6_L 
generic map(
  INIT => X"FFFFFFFFFFFFFFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1711\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1648\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1710\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_2_0\(17),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1661\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_1\(17),
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_REP2\(17));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2_Z8596\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP2\,
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_REP2\(17),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIIH1P3[230]\: LUT6 
generic map(
  INIT => X"135FECA00000FFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(230),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_1_N_4_3\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_1_N_6_7\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST_RNIKBRQ1[8]\: LUT5_L 
generic map(
  INIT => X"070F77FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_FAST\(8),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(11),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_1_N_6_7\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS_2_RNIVG5P[1]\: LUT4 
generic map(
  INIT => X"B847"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(114),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_17_REP1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS_2\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_AXB_1_N_4_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_FAST[9]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7908\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7732\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7968\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_FAST\(9));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_REP1[9]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7908\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7732\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7968\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_REP1\(9));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_FAST[7]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7910\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7734\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7970\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_FAST\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_REP1[7]\: LUT5_L 
generic map(
  INIT => X"FEBA5410"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7910\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7734\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7970\,
  LO => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_REP1\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_I_155\: MUXCY port map (
    DI => NN_2,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_DATA_TMP\(18),
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_0_N_3_I\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_I_35\: MUXCY port map (
    DI => NN_2,
    CI => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_0_DATA_TMP\(3),
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12030\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS\);
\GRLFPC20.R.X.RDD_GRLFPC20.R.X.SEQERR_1\: SRL16E port map (
  Q => \GRLFPC20.R.X.RDD_TMP_D_ARRAY_0\(0),
  A0 => NN_2,
  A1 => NN_3,
  A2 => NN_2,
  A3 => NN_2,
  D => \GRLFPC20.COMB.RDD_1\,
  CLK => clk,
  CE => holdn);
\GRLFPC20.R.X.SEQERR_GRLFPC20.R.X.SEQERR_1\: SRL16E port map (
  Q => \GRLFPC20.R.X.SEQERR_TMP_D_ARRAY_0\(0),
  A0 => NN_2,
  A1 => NN_3,
  A2 => NN_2,
  A3 => NN_2,
  D => \GRLFPC20.COMB.V.A.SEQERR_1\,
  CLK => clk,
  CE => holdn);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_7_REP1_Z8608\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_7_REP1\,
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_REP1\(7),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST[7]_Z8609\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST\(7),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_FAST\(7),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_9_REP1_Z8610\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_9_REP1\,
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_REP1\(9),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST[9]_Z8611\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST\(9),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_FAST\(9),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_8_REP1_Z8612\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_8_REP1\,
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_REP1\(8),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST[8]_Z8613\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST\(8),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_FAST\(8),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2_Z8614\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_10\(10),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1_Z8615\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1\,
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_10\(10),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_FAST[10]_Z8616\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_FAST\(10),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_10\(10),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST[17]_Z8617\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST\(17),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_FAST\(17),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST[15]_Z8618\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST\(15),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_FAST\(15),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_3_REP1_Z8619\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_3_REP1\,
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_REP1\(3),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST[3]_Z8620\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST\(3),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_FAST\(3),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST[376]_Z8621\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST\(376),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_DIVMULTV_FAST\(0),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST[1]_Z8622\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST\(1),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1_FAST\(1),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST[374]_Z8623\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_FAST\(374),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_FAST\(374),
    C => clk);
\GRLFPC20.R.X.RDD_DOUT[0]\: FDE port map (
    Q => \GRLFPC20.R.X.RDD\,
    D => \GRLFPC20.R.X.RDD_TMP_D_ARRAY_0\(0),
    C => clk,
    CE => holdn);
\GRLFPC20.R.X.SEQERR_DOUT[0]\: FDE port map (
    Q => \GRLFPC20.R.X.SEQERR\,
    D => \GRLFPC20.R.X.SEQERR_TMP_D_ARRAY_0\(0),
    C => clk,
    CE => holdn);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RET_Z8626\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RET\,
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8537_RETI\,
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.R.MK.HOLDN2_Z8627\: FD port map (
    Q => \GRLFPC20.R.MK.HOLDN2\,
    D => \GRLFPC20.R.MK.HOLDN1\,
    C => clk);
\GRLFPC20.R.MK.RST2_Z8628\: FD port map (
    Q => \GRLFPC20.R.MK.RST2\,
    D => \GRLFPC20.R.MK.RST\,
    C => clk);
\GRLFPC20.R.MK.RST_Z8629\: FD port map (
    Q => \GRLFPC20.R.MK.RST\,
    D => \GRLFPC20.COMB.V.MK.RST_1\,
    C => clk);
\GRLFPC20.R.A.RS1[0]_Z8630\: FD port map (
    Q => \GRLFPC20.R.A.RS1\(0),
    D => \GRLFPC20.COMB.RS1_1\(0),
    C => clk);
\GRLFPC20.R.I.RES[7]_Z8631\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(7),
    D => \GRLFPC20.FPO.FRAC\(10),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[6]_Z8632\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(6),
    D => \GRLFPC20.FPO.FRAC\(9),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[5]_Z8633\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(5),
    D => \GRLFPC20.FPO.FRAC\(8),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[4]_Z8634\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(4),
    D => \GRLFPC20.FPO.FRAC\(7),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[3]_Z8635\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(3),
    D => \GRLFPC20.FPO.FRAC\(6),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[2]_Z8636\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(2),
    D => \GRLFPC20.FPO.FRAC\(5),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[1]_Z8637\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(1),
    D => \GRLFPC20.FPO.FRAC\(4),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[0]_Z8638\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(0),
    D => \GRLFPC20.FPO.FRAC\(3),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[22]_Z8639\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(22),
    D => \GRLFPC20.FPO.FRAC\(25),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[21]_Z8640\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(21),
    D => \GRLFPC20.FPO.FRAC\(24),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[20]_Z8641\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(20),
    D => \GRLFPC20.FPO.FRAC\(23),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[19]_Z8642\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(19),
    D => \GRLFPC20.FPO.FRAC\(22),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[18]_Z8643\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(18),
    D => \GRLFPC20.FPO.FRAC\(21),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[17]_Z8644\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(17),
    D => \GRLFPC20.FPO.FRAC\(20),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[16]_Z8645\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(16),
    D => \GRLFPC20.FPO.FRAC\(19),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[15]_Z8646\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(15),
    D => \GRLFPC20.FPO.FRAC\(18),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[14]_Z8647\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(14),
    D => \GRLFPC20.FPO.FRAC\(17),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[13]_Z8648\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(13),
    D => \GRLFPC20.FPO.FRAC\(16),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[12]_Z8649\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(12),
    D => \GRLFPC20.FPO.FRAC\(15),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[11]_Z8650\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(11),
    D => \GRLFPC20.FPO.FRAC\(14),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[10]_Z8651\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(10),
    D => \GRLFPC20.FPO.FRAC\(13),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[9]_Z8652\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(9),
    D => \GRLFPC20.FPO.FRAC\(12),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[8]_Z8653\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(8),
    D => \GRLFPC20.FPO.FRAC\(11),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[37]_Z8654\: FD port map (
    Q => \GRLFPC20.R.I.RES\(37),
    D => \GRLFPC20.COMB.V.I.RES_1\(37),
    C => clk);
\GRLFPC20.R.I.RES[36]_Z8655\: FD port map (
    Q => \GRLFPC20.R.I.RES\(36),
    D => \GRLFPC20.COMB.V.I.RES_1\(36),
    C => clk);
\GRLFPC20.R.I.RES[35]_Z8656\: FD port map (
    Q => \GRLFPC20.R.I.RES\(35),
    D => \GRLFPC20.COMB.V.I.RES_1\(35),
    C => clk);
\GRLFPC20.R.I.RES[34]_Z8657\: FD port map (
    Q => \GRLFPC20.R.I.RES\(34),
    D => \GRLFPC20.COMB.V.I.RES_1\(34),
    C => clk);
\GRLFPC20.R.I.RES[33]_Z8658\: FD port map (
    Q => \GRLFPC20.R.I.RES\(33),
    D => \GRLFPC20.COMB.V.I.RES_1\(33),
    C => clk);
\GRLFPC20.R.I.RES[32]_Z8659\: FD port map (
    Q => \GRLFPC20.R.I.RES\(32),
    D => \GRLFPC20.COMB.V.I.RES_1\(32),
    C => clk);
\GRLFPC20.R.I.RES[31]_Z8660\: FD port map (
    Q => \GRLFPC20.R.I.RES\(31),
    D => \GRLFPC20.COMB.V.I.RES_1\(31),
    C => clk);
\GRLFPC20.R.I.RES[30]_Z8661\: FD port map (
    Q => \GRLFPC20.R.I.RES\(30),
    D => \GRLFPC20.COMB.V.I.RES_1\(30),
    C => clk);
\GRLFPC20.R.I.RES[29]_Z8662\: FD port map (
    Q => \GRLFPC20.R.I.RES\(29),
    D => \GRLFPC20.COMB.V.I.RES_1\(29),
    C => clk);
\GRLFPC20.R.I.RES[28]_Z8663\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(28),
    D => \GRLFPC20.FPO.FRAC\(31),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[27]_Z8664\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(27),
    D => \GRLFPC20.FPO.FRAC\(30),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[26]_Z8665\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(26),
    D => \GRLFPC20.FPO.FRAC\(29),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[25]_Z8666\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(25),
    D => \GRLFPC20.FPO.FRAC\(28),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[24]_Z8667\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(24),
    D => \GRLFPC20.FPO.FRAC\(27),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[23]_Z8668\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(23),
    D => \GRLFPC20.FPO.FRAC\(26),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[52]_Z8669\: FD port map (
    Q => \GRLFPC20.R.I.RES\(52),
    D => \GRLFPC20.COMB.V.I.RES_1\(52),
    C => clk);
\GRLFPC20.R.I.RES[51]_Z8670\: FD port map (
    Q => \GRLFPC20.R.I.RES\(51),
    D => \GRLFPC20.COMB.V.I.RES_1\(51),
    C => clk);
\GRLFPC20.R.I.RES[50]_Z8671\: FD port map (
    Q => \GRLFPC20.R.I.RES\(50),
    D => \GRLFPC20.COMB.V.I.RES_1\(50),
    C => clk);
\GRLFPC20.R.I.RES[49]_Z8672\: FD port map (
    Q => \GRLFPC20.R.I.RES\(49),
    D => \GRLFPC20.COMB.V.I.RES_1\(49),
    C => clk);
\GRLFPC20.R.I.RES[48]_Z8673\: FD port map (
    Q => \GRLFPC20.R.I.RES\(48),
    D => \GRLFPC20.COMB.V.I.RES_1\(48),
    C => clk);
\GRLFPC20.R.I.RES[47]_Z8674\: FD port map (
    Q => \GRLFPC20.R.I.RES\(47),
    D => \GRLFPC20.COMB.V.I.RES_1\(47),
    C => clk);
\GRLFPC20.R.I.RES[46]_Z8675\: FD port map (
    Q => \GRLFPC20.R.I.RES\(46),
    D => \GRLFPC20.COMB.V.I.RES_1\(46),
    C => clk);
\GRLFPC20.R.I.RES[45]_Z8676\: FD port map (
    Q => \GRLFPC20.R.I.RES\(45),
    D => \GRLFPC20.COMB.V.I.RES_1\(45),
    C => clk);
\GRLFPC20.R.I.RES[44]_Z8677\: FD port map (
    Q => \GRLFPC20.R.I.RES\(44),
    D => \GRLFPC20.COMB.V.I.RES_1\(44),
    C => clk);
\GRLFPC20.R.I.RES[43]_Z8678\: FD port map (
    Q => \GRLFPC20.R.I.RES\(43),
    D => \GRLFPC20.COMB.V.I.RES_1\(43),
    C => clk);
\GRLFPC20.R.I.RES[42]_Z8679\: FD port map (
    Q => \GRLFPC20.R.I.RES\(42),
    D => \GRLFPC20.COMB.V.I.RES_1\(42),
    C => clk);
\GRLFPC20.R.I.RES[41]_Z8680\: FD port map (
    Q => \GRLFPC20.R.I.RES\(41),
    D => \GRLFPC20.COMB.V.I.RES_1\(41),
    C => clk);
\GRLFPC20.R.I.RES[40]_Z8681\: FD port map (
    Q => \GRLFPC20.R.I.RES\(40),
    D => \GRLFPC20.COMB.V.I.RES_1\(40),
    C => clk);
\GRLFPC20.R.I.RES[39]_Z8682\: FD port map (
    Q => \GRLFPC20.R.I.RES\(39),
    D => \GRLFPC20.COMB.V.I.RES_1\(39),
    C => clk);
\GRLFPC20.R.I.RES[38]_Z8683\: FD port map (
    Q => \GRLFPC20.R.I.RES\(38),
    D => \GRLFPC20.COMB.V.I.RES_1\(38),
    C => clk);
\GRLFPC20.R.I.RES[63]_Z8684\: FD port map (
    Q => \GRLFPC20.R.I.RES\(63),
    D => \GRLFPC20.COMB.V.I.RES_1\(63),
    C => clk);
\GRLFPC20.R.I.RES[62]_Z8685\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(62),
    D => \GRLFPC20.FPO.EXP\(10),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[61]_Z8686\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(61),
    D => \GRLFPC20.FPO.EXP\(9),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[60]_Z8687\: FDE port map (
    Q => \GRLFPC20.R.I.RES\(60),
    D => \GRLFPC20.FPO.EXP\(8),
    C => clk,
    CE => \GRLFPC20.N_2102\);
\GRLFPC20.R.I.RES[59]_Z8688\: FD port map (
    Q => \GRLFPC20.R.I.RES\(59),
    D => \GRLFPC20.COMB.V.I.RES_1\(59),
    C => clk);
\GRLFPC20.R.I.RES[58]_Z8689\: FD port map (
    Q => \GRLFPC20.R.I.RES\(58),
    D => \GRLFPC20.COMB.V.I.RES_1\(58),
    C => clk);
\GRLFPC20.R.I.RES[57]_Z8690\: FD port map (
    Q => \GRLFPC20.R.I.RES\(57),
    D => \GRLFPC20.COMB.V.I.RES_1\(57),
    C => clk);
\GRLFPC20.R.I.RES[56]_Z8691\: FD port map (
    Q => \GRLFPC20.R.I.RES\(56),
    D => \GRLFPC20.COMB.V.I.RES_1\(56),
    C => clk);
\GRLFPC20.R.I.RES[55]_Z8692\: FD port map (
    Q => \GRLFPC20.R.I.RES\(55),
    D => \GRLFPC20.COMB.V.I.RES_1\(55),
    C => clk);
\GRLFPC20.R.I.RES[54]_Z8693\: FD port map (
    Q => \GRLFPC20.R.I.RES\(54),
    D => \GRLFPC20.COMB.V.I.RES_1\(54),
    C => clk);
\GRLFPC20.R.I.RES[53]_Z8694\: FD port map (
    Q => \GRLFPC20.R.I.RES\(53),
    D => \GRLFPC20.COMB.V.I.RES_1\(53),
    C => clk);
\GRLFPC20.R.E.AFQ_Z8695\: FDE port map (
    Q => \GRLFPC20.R.E.AFQ\,
    D => \GRLFPC20.COMB.V.E.AFQ_1\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.AFSR_Z8696\: FDE port map (
    Q => \GRLFPC20.R.E.AFSR\,
    D => \GRLFPC20.COMB.V.E.AFSR_1\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.FPOP_Z8697\: FDE port map (
    Q => \GRLFPC20.R.E.FPOP\,
    D => \GRLFPC20.N_2931_1\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.LD_Z8698\: FDE port map (
    Q => \GRLFPC20.R.E.LD\,
    D => \GRLFPC20.COMB.V.E.LD_1\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.M.AFQ_Z8699\: FDE port map (
    Q => \GRLFPC20.R.M.AFQ\,
    D => \GRLFPC20.COMB.V.M.AFQ_1\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.M.AFSR_Z8700\: FDE port map (
    Q => \GRLFPC20.R.M.AFSR\,
    D => \GRLFPC20.COMB.V.M.AFSR_1\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.M.FPOP_Z8701\: FDE port map (
    Q => \GRLFPC20.R.M.FPOP\,
    D => \GRLFPC20.COMB.V.M.FPOP_1\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.M.LD_Z8702\: FDE port map (
    Q => \GRLFPC20.R.M.LD\,
    D => \GRLFPC20.COMB.V.M.LD_1\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.X.AFQ_Z8703\: FDE port map (
    Q => \GRLFPC20.R.X.AFQ\,
    D => \GRLFPC20.COMB.V.X.AFQ_1\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.X.AFSR_Z8704\: FDE port map (
    Q => \GRLFPC20.R.X.AFSR\,
    D => \GRLFPC20.COMB.V.X.AFSR_1\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.X.FPOP_Z8705\: FDE port map (
    Q => \GRLFPC20.R.X.FPOP\,
    D => \GRLFPC20.COMB.V.X.FPOP_1\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.X.LD_Z8706\: FDE port map (
    Q => \GRLFPC20.R.X.LD\,
    D => \GRLFPC20.COMB.V.X.LD_1\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.I.PC[31]_Z8707\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(31),
    D => cpi_x_pc(31),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[30]_Z8708\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(30),
    D => cpi_x_pc(30),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[29]_Z8709\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(29),
    D => cpi_x_pc(29),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[28]_Z8710\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(28),
    D => cpi_x_pc(28),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[27]_Z8711\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(27),
    D => cpi_x_pc(27),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[26]_Z8712\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(26),
    D => cpi_x_pc(26),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[25]_Z8713\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(25),
    D => cpi_x_pc(25),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[24]_Z8714\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(24),
    D => cpi_x_pc(24),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[23]_Z8715\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(23),
    D => cpi_x_pc(23),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[22]_Z8716\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(22),
    D => cpi_x_pc(22),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[21]_Z8717\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(21),
    D => cpi_x_pc(21),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[20]_Z8718\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(20),
    D => cpi_x_pc(20),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[19]_Z8719\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(19),
    D => cpi_x_pc(19),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[18]_Z8720\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(18),
    D => cpi_x_pc(18),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[17]_Z8721\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(17),
    D => cpi_x_pc(17),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[16]_Z8722\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(16),
    D => cpi_x_pc(16),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[15]_Z8723\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(15),
    D => cpi_x_pc(15),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[14]_Z8724\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(14),
    D => cpi_x_pc(14),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[13]_Z8725\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(13),
    D => cpi_x_pc(13),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[12]_Z8726\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(12),
    D => cpi_x_pc(12),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[11]_Z8727\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(11),
    D => cpi_x_pc(11),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[10]_Z8728\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(10),
    D => cpi_x_pc(10),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[9]_Z8729\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(9),
    D => cpi_x_pc(9),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[8]_Z8730\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(8),
    D => cpi_x_pc(8),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[7]_Z8731\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(7),
    D => cpi_x_pc(7),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[6]_Z8732\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(6),
    D => cpi_x_pc(6),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[5]_Z8733\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(5),
    D => cpi_x_pc(5),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[4]_Z8734\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(4),
    D => cpi_x_pc(4),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[3]_Z8735\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(3),
    D => cpi_x_pc(3),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.I.PC[2]_Z8736\: FDE port map (
    Q => \GRLFPC20.R.I.PC\(2),
    D => cpi_x_pc(2),
    C => clk,
    CE => N_3710);
\GRLFPC20.R.A.MOV_Z8737\: FDE port map (
    Q => \GRLFPC20.R.A.MOV\,
    D => \GRLFPC20.N_865\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.I.RDD_Z8738\: FDE port map (
    Q => \GRLFPC20.R.I.RDD\,
    D => \GRLFPC20.N_3022_I\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[31]\: FDE port map (
    Q => cpo_data(31),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(31),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[30]\: FDE port map (
    Q => cpo_data(30),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(30),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[29]\: FDE port map (
    Q => cpo_data(29),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(29),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[28]\: FDE port map (
    Q => cpo_data(28),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(28),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[27]\: FDE port map (
    Q => cpo_data(27),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(27),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[26]\: FDE port map (
    Q => cpo_data(26),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(26),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[25]\: FDE port map (
    Q => cpo_data(25),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(25),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[24]\: FDE port map (
    Q => cpo_data(24),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(24),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[23]\: FDE port map (
    Q => cpo_data(23),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(23),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[22]\: FDE port map (
    Q => cpo_data(22),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(22),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[21]\: FDE port map (
    Q => cpo_data(21),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(21),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[20]\: FDE port map (
    Q => cpo_data(20),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(20),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[19]\: FDE port map (
    Q => cpo_data(19),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(19),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[18]\: FDE port map (
    Q => cpo_data(18),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(18),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[17]\: FDE port map (
    Q => cpo_data(17),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(17),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[16]\: FDE port map (
    Q => cpo_data(16),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(16),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[15]\: FDE port map (
    Q => cpo_data(15),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(15),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[14]\: FDE port map (
    Q => cpo_data(14),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(14),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[13]\: FDE port map (
    Q => cpo_data(13),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(13),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[12]\: FDE port map (
    Q => cpo_data(12),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(12),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[11]\: FDE port map (
    Q => cpo_data(11),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(11),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[10]\: FDE port map (
    Q => cpo_data(10),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(10),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[9]\: FDE port map (
    Q => cpo_data(9),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(9),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[8]\: FDE port map (
    Q => cpo_data(8),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(8),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[7]\: FDE port map (
    Q => cpo_data(7),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(7),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[6]\: FDE port map (
    Q => cpo_data(6),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(6),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[5]\: FDE port map (
    Q => cpo_data(5),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(5),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[4]\: FDE port map (
    Q => cpo_data(4),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(4),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[3]\: FDE port map (
    Q => cpo_data(3),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(3),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[2]\: FDE port map (
    Q => cpo_data(2),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(2),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[1]\: FDE port map (
    Q => cpo_data(1),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(1),
    C => clk,
    CE => holdn);
\GRLFPC20.R.E.STDATA[0]\: FDE port map (
    Q => cpo_data(0),
    D => \GRLFPC20.COMB.V.E.STDATA_1\(0),
    C => clk,
    CE => holdn);
\GRLFPC20.R.FSR.NONSTD_Z8771\: FDE port map (
    Q => \GRLFPC20.R.FSR.NONSTD\,
    D => \GRLFPC20.COMB.V.FSR.NONSTD_1\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.FSR.RD[1]_Z8772\: FDE port map (
    Q => \GRLFPC20.R.FSR.RD\(1),
    D => \GRLFPC20.COMB.V.FSR.RD_1\(1),
    C => clk,
    CE => holdn);
\GRLFPC20.R.FSR.RD[0]_Z8773\: FDE port map (
    Q => \GRLFPC20.R.FSR.RD\(0),
    D => \GRLFPC20.COMB.V.FSR.RD_1\(0),
    C => clk,
    CE => holdn);
\GRLFPC20.R.FSR.TEM[4]_Z8774\: FDE port map (
    Q => \GRLFPC20.R.FSR.TEM\(4),
    D => \GRLFPC20.COMB.V.FSR.TEM_1\(4),
    C => clk,
    CE => holdn);
\GRLFPC20.R.FSR.TEM[3]_Z8775\: FDE port map (
    Q => \GRLFPC20.R.FSR.TEM\(3),
    D => \GRLFPC20.COMB.V.FSR.TEM_1\(3),
    C => clk,
    CE => holdn);
\GRLFPC20.R.FSR.TEM[2]_Z8776\: FDE port map (
    Q => \GRLFPC20.R.FSR.TEM\(2),
    D => \GRLFPC20.COMB.V.FSR.TEM_1\(2),
    C => clk,
    CE => holdn);
\GRLFPC20.R.FSR.TEM[1]_Z8777\: FDE port map (
    Q => \GRLFPC20.R.FSR.TEM\(1),
    D => \GRLFPC20.COMB.V.FSR.TEM_1\(1),
    C => clk,
    CE => holdn);
\GRLFPC20.R.FSR.TEM[0]_Z8778\: FDE port map (
    Q => \GRLFPC20.R.FSR.TEM\(0),
    D => \GRLFPC20.COMB.V.FSR.TEM_1\(0),
    C => clk,
    CE => holdn);
\GRLFPC20.R.A.RS2D_Z8779\: FDE port map (
    Q => \GRLFPC20.R.A.RS2D\,
    D => \GRLFPC20.COMB.RS2D_1\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.A.RS1D_Z8780\: FDE port map (
    Q => \GRLFPC20.R.A.RS1D\,
    D => \GRLFPC20.COMB.RS1D_1\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.STATE[1]_Z8781\: FDE port map (
    Q => \GRLFPC20.R.STATE\(1),
    D => \GRLFPC20.COMB.V.STATE_1_IV_I\(1),
    C => clk,
    CE => holdn);
\GRLFPC20.R.STATE[0]_Z8782\: FDE port map (
    Q => \GRLFPC20.R.STATE\(0),
    D => \GRLFPC20.COMB.V.STATE_1\(0),
    C => clk,
    CE => holdn);
\GRLFPC20.R.FSR.FTT[2]_Z8783\: FDE port map (
    Q => \GRLFPC20.R.FSR.FTT\(2),
    D => \GRLFPC20.COMB.V.FSR.FTT_1\(2),
    C => clk,
    CE => holdn);
\GRLFPC20.R.FSR.FTT[1]_Z8784\: FDE port map (
    Q => \GRLFPC20.R.FSR.FTT\(1),
    D => \GRLFPC20.COMB.V.FSR.FTT_1\(1),
    C => clk,
    CE => holdn);
\GRLFPC20.R.FSR.FTT[0]_Z8785\: FDE port map (
    Q => \GRLFPC20.R.FSR.FTT\(0),
    D => \GRLFPC20.COMB.V.FSR.FTT_1\(0),
    C => clk,
    CE => holdn);
\GRLFPC20.R.A.RF2REN[1]_Z8786\: FDE port map (
    Q => \GRLFPC20.R.A.RF2REN\(1),
    D => \GRLFPC20.N_2961_I\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.A.RF2REN[2]_Z8787\: FDE port map (
    Q => \GRLFPC20.R.A.RF2REN\(2),
    D => \GRLFPC20.N_2941_I\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.A.AFQ_Z8788\: FDE port map (
    Q => \GRLFPC20.R.A.AFQ\,
    D => \GRLFPC20.COMB.V.A.AFQ_1\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.A.AFSR_Z8789\: FDE port map (
    Q => \GRLFPC20.R.A.AFSR\,
    D => \GRLFPC20.COMB.V.A.AFSR_1\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.A.FPOP_Z8790\: FDE port map (
    Q => \GRLFPC20.R.A.FPOP\,
    D => \GRLFPC20.N_1312\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.A.LD_Z8791\: FDE port map (
    Q => \GRLFPC20.R.A.LD\,
    D => \GRLFPC20.COMB.V.A.LD_1\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.A.ST_Z8792\: FDE port map (
    Q => \GRLFPC20.R.A.ST\,
    D => \GRLFPC20.COMB.V.A.ST_1\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.I.EXEC_Z8793\: FDE port map (
    Q => \GRLFPC20.R.I.EXEC\,
    D => \GRLFPC20.N_2929_I\,
    C => clk,
    CE => holdn);
\GRLFPC20.R.FSR.FCC[1]\: FDE port map (
    Q => CPO_CC_3,
    D => \GRLFPC20.COMB.V.FSR.FCC_1\(1),
    C => clk,
    CE => holdn);
\GRLFPC20.R.FSR.FCC[0]\: FDE port map (
    Q => NN_1,
    D => \GRLFPC20.COMB.V.FSR.FCC_1\(0),
    C => clk,
    CE => holdn);
\GRLFPC20.R.FSR.AEXC[4]_Z8796\: FDE port map (
    Q => \GRLFPC20.R.FSR.AEXC\(4),
    D => \GRLFPC20.COMB.V.FSR.AEXC_1\(4),
    C => clk,
    CE => holdn);
\GRLFPC20.R.FSR.AEXC[3]_Z8797\: FDE port map (
    Q => \GRLFPC20.R.FSR.AEXC\(3),
    D => \GRLFPC20.COMB.V.FSR.AEXC_1\(3),
    C => clk,
    CE => holdn);
\GRLFPC20.R.FSR.AEXC[2]_Z8798\: FDE port map (
    Q => \GRLFPC20.R.FSR.AEXC\(2),
    D => \GRLFPC20.COMB.V.FSR.AEXC_1\(2),
    C => clk,
    CE => holdn);
\GRLFPC20.R.FSR.AEXC[1]_Z8799\: FDE port map (
    Q => \GRLFPC20.R.FSR.AEXC\(1),
    D => \GRLFPC20.COMB.V.FSR.AEXC_1\(1),
    C => clk,
    CE => holdn);
\GRLFPC20.R.FSR.AEXC[0]_Z8800\: FDE port map (
    Q => \GRLFPC20.R.FSR.AEXC\(0),
    D => \GRLFPC20.COMB.V.FSR.AEXC_1\(0),
    C => clk,
    CE => holdn);
\GRLFPC20.R.FSR.CEXC[4]_Z8801\: FDE port map (
    Q => \GRLFPC20.R.FSR.CEXC\(4),
    D => \GRLFPC20.COMB.V.FSR.CEXC_1\(4),
    C => clk,
    CE => holdn);
\GRLFPC20.R.FSR.CEXC[3]_Z8802\: FDE port map (
    Q => \GRLFPC20.R.FSR.CEXC\(3),
    D => \GRLFPC20.COMB.V.FSR.CEXC_1\(3),
    C => clk,
    CE => holdn);
\GRLFPC20.R.FSR.CEXC[2]_Z8803\: FDE port map (
    Q => \GRLFPC20.R.FSR.CEXC\(2),
    D => \GRLFPC20.COMB.V.FSR.CEXC_1\(2),
    C => clk,
    CE => holdn);
\GRLFPC20.R.FSR.CEXC[1]_Z8804\: FDE port map (
    Q => \GRLFPC20.R.FSR.CEXC\(1),
    D => \GRLFPC20.COMB.V.FSR.CEXC_1\(1),
    C => clk,
    CE => holdn);
\GRLFPC20.R.FSR.CEXC[0]_Z8805\: FDE port map (
    Q => \GRLFPC20.R.FSR.CEXC\(0),
    D => \GRLFPC20.COMB.V.FSR.CEXC_1\(0),
    C => clk,
    CE => holdn);
\GRLFPC20.R.I.V_Z8806\: FDR port map (
    Q => \GRLFPC20.R.I.V\,
    D => \GRLFPC20.R.I.V_0\,
    C => clk,
    R => RST_I);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL[4]_Z8807\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(4),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_14\(4),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL[7]_Z8808\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(7),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL[10]_Z8809\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_10\(10),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL[11]_Z8810\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
    D => CPI_D_INST_I(6),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL[12]_Z8811\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(12),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9260\,
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL[13]_Z8812\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(13),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9252\,
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL[14]_Z8813\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(14),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_871_I\,
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL[15]_Z8814\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(42),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL[16]_Z8815\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(16),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_870_I\,
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL[3]_Z8816\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(3),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_13\(3),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[376]_Z8817\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(376),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_DIVMULTV\(0),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[377]_Z8818\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(377),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_I\(0),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[361]_Z8819\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(361),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(102),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[362]_Z8820\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(362),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(103),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[363]_Z8821\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(363),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(104),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[364]_Z8822\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(364),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(105),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[365]_Z8823\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(365),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(106),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[366]_Z8824\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(366),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(107),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[367]_Z8825\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(367),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(108),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[368]_Z8826\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(368),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(109),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[369]_Z8827\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(369),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(110),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[370]_Z8828\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(370),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(111),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[371]_Z8829\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(371),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(112),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[372]_Z8830\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(372),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(113),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[373]_Z8831\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(373),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_25_I\(0),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[374]_Z8832\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(374),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(374),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[375]_Z8833\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(375),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(375),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[346]_Z8834\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(346),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(87),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[347]_Z8835\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(347),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(88),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[348]_Z8836\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(348),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(89),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[349]_Z8837\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(349),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(90),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[350]_Z8838\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(350),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(91),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[351]_Z8839\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(351),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(92),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[352]_Z8840\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(352),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(93),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[353]_Z8841\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(353),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(94),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[354]_Z8842\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(354),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(95),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[355]_Z8843\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(355),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(96),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[356]_Z8844\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(356),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(97),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[357]_Z8845\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(357),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(98),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[358]_Z8846\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(358),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(99),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[359]_Z8847\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(359),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(100),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[360]_Z8848\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(360),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(101),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[331]_Z8849\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(331),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(72),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[332]_Z8850\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(332),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(73),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[333]_Z8851\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(333),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(74),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[334]_Z8852\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(334),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(75),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[335]_Z8853\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(335),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(76),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[336]_Z8854\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(336),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(77),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[337]_Z8855\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(337),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(78),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[338]_Z8856\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(338),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(79),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[339]_Z8857\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(339),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(80),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[340]_Z8858\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(340),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(81),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[341]_Z8859\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(341),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(82),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[342]_Z8860\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(342),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(83),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[343]_Z8861\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(343),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(84),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[344]_Z8862\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(344),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(85),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[345]_Z8863\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(345),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(86),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[316]_Z8864\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(316),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_50\(316),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[317]_Z8865\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(317),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(58),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[318]_Z8866\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(318),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(59),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[319]_Z8867\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(319),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(60),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[320]_Z8868\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(320),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(61),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[321]_Z8869\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(321),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(62),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[322]_Z8870\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(322),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(63),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[323]_Z8871\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(323),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(64),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[324]_Z8872\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(324),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(65),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[325]_Z8873\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(325),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(66),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[326]_Z8874\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(326),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(67),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[327]_Z8875\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(327),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(68),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[328]_Z8876\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(328),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(69),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[329]_Z8877\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(329),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(70),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[330]_Z8878\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(330),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(71),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[301]_Z8879\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(301),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(42),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[302]_Z8880\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(302),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(43),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[303]_Z8881\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(303),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(44),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[304]_Z8882\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(304),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(45),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[305]_Z8883\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(305),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(46),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[306]_Z8884\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(306),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(47),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[307]_Z8885\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(307),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(48),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[308]_Z8886\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(308),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(49),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[309]_Z8887\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(309),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(50),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[310]_Z8888\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(310),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(51),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[311]_Z8889\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(311),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(52),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[312]_Z8890\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(312),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(53),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[313]_Z8891\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(313),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(54),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[314]_Z8892\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(314),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(55),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[315]_Z8893\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(315),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(57),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[286]_Z8894\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(286),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(27),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[287]_Z8895\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(287),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(28),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[288]_Z8896\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(288),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(29),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[289]_Z8897\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(289),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(30),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[290]_Z8898\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(290),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(31),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[291]_Z8899\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(291),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(32),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[292]_Z8900\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(292),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(33),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[293]_Z8901\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(293),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(34),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[294]_Z8902\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(294),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(35),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[295]_Z8903\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(295),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(36),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[296]_Z8904\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(296),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(37),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[297]_Z8905\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(297),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(38),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[298]_Z8906\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(298),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(39),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[299]_Z8907\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(299),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(40),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[300]_Z8908\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(300),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(41),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[271]_Z8909\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(271),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(12),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[272]_Z8910\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(272),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(13),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[273]_Z8911\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(273),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(14),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[274]_Z8912\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(274),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(15),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[275]_Z8913\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(275),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(16),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[276]_Z8914\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(276),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(17),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[277]_Z8915\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(277),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(18),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[278]_Z8916\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(278),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(19),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[279]_Z8917\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(279),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(20),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[280]_Z8918\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(280),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(21),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[281]_Z8919\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(281),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(22),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[282]_Z8920\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(282),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(23),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[283]_Z8921\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(283),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(24),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[284]_Z8922\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(284),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(25),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[285]_Z8923\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(285),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(26),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[258]_Z8924\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(258),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_49\(258),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[259]_Z8925\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(259),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(0),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[260]_Z8926\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(260),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(1),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[261]_Z8927\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(261),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(2),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[262]_Z8928\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(262),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12045_I\,
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[263]_Z8929\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(263),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(4),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[264]_Z8930\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(264),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(5),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[265]_Z8931\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(265),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(6),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[266]_Z8932\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(266),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(7),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[267]_Z8933\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(267),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(8),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[268]_Z8934\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(268),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(9),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[269]_Z8935\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(269),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(10),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[270]_Z8936\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(270),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(11),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[241]_Z8937\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(241),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(241),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[242]_Z8938\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(242),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(242),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[243]_Z8939\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(243),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(243),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[244]_Z8940\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(244),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[247]_Z8941\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(247),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(247),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[248]_Z8942\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(248),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(248),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[249]_Z8943\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(249),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(249),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[226]_Z8944\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(226),
    D => \GRLFPC20.FPO.FRAC\(5),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[227]_Z8945\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(227),
    D => \GRLFPC20.FPO.FRAC\(4),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[228]_Z8946\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(228),
    D => \GRLFPC20.FPO.FRAC\(3),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[229]_Z8947\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(229),
    D => N_3827,
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[230]_Z8948\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(230),
    D => N_3826,
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[231]_Z8949\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(231),
    D => N_3825,
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[237]_Z8950\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(237),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(237),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[238]_Z8951\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(238),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(238),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[239]_Z8952\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(239),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(239),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[240]_Z8953\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(240),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(240),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[211]_Z8954\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(211),
    D => \GRLFPC20.FPO.FRAC\(20),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[212]_Z8955\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(212),
    D => \GRLFPC20.FPO.FRAC\(19),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[213]_Z8956\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(213),
    D => \GRLFPC20.FPO.FRAC\(18),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[214]_Z8957\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(214),
    D => \GRLFPC20.FPO.FRAC\(17),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[215]_Z8958\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(215),
    D => \GRLFPC20.FPO.FRAC\(16),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[216]_Z8959\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(216),
    D => \GRLFPC20.FPO.FRAC\(15),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[217]_Z8960\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(217),
    D => \GRLFPC20.FPO.FRAC\(14),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[218]_Z8961\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(218),
    D => \GRLFPC20.FPO.FRAC\(13),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[219]_Z8962\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(219),
    D => \GRLFPC20.FPO.FRAC\(12),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[220]_Z8963\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(220),
    D => \GRLFPC20.FPO.FRAC\(11),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[221]_Z8964\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(221),
    D => \GRLFPC20.FPO.FRAC\(10),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[222]_Z8965\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(222),
    D => \GRLFPC20.FPO.FRAC\(9),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[223]_Z8966\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(223),
    D => \GRLFPC20.FPO.FRAC\(8),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[224]_Z8967\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(224),
    D => \GRLFPC20.FPO.FRAC\(7),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[225]_Z8968\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(225),
    D => \GRLFPC20.FPO.FRAC\(6),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[196]_Z8969\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(196),
    D => \GRLFPC20.FPO.FRAC\(35),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[197]_Z8970\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(197),
    D => \GRLFPC20.FPO.FRAC\(34),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[198]_Z8971\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(198),
    D => \GRLFPC20.FPO.FRAC\(33),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[199]_Z8972\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(199),
    D => \GRLFPC20.FPO.FRAC\(32),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[200]_Z8973\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(200),
    D => \GRLFPC20.FPO.FRAC\(31),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[201]_Z8974\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(201),
    D => \GRLFPC20.FPO.FRAC\(30),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[202]_Z8975\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(202),
    D => \GRLFPC20.FPO.FRAC\(29),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[203]_Z8976\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(203),
    D => \GRLFPC20.FPO.FRAC\(28),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[204]_Z8977\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(204),
    D => \GRLFPC20.FPO.FRAC\(27),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[205]_Z8978\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(205),
    D => \GRLFPC20.FPO.FRAC\(26),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[206]_Z8979\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(206),
    D => \GRLFPC20.FPO.FRAC\(25),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[207]_Z8980\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(207),
    D => \GRLFPC20.FPO.FRAC\(24),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[208]_Z8981\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(208),
    D => \GRLFPC20.FPO.FRAC\(23),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[209]_Z8982\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(209),
    D => \GRLFPC20.FPO.FRAC\(22),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[210]_Z8983\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(210),
    D => \GRLFPC20.FPO.FRAC\(21),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[181]_Z8984\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(181),
    D => \GRLFPC20.FPO.FRAC\(50),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[182]_Z8985\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(182),
    D => \GRLFPC20.FPO.FRAC\(49),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[183]_Z8986\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(183),
    D => \GRLFPC20.FPO.FRAC\(48),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[184]_Z8987\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(184),
    D => \GRLFPC20.FPO.FRAC\(47),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[185]_Z8988\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(185),
    D => \GRLFPC20.FPO.FRAC\(46),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[186]_Z8989\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(186),
    D => \GRLFPC20.FPO.FRAC\(45),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[187]_Z8990\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(187),
    D => \GRLFPC20.FPO.FRAC\(44),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[188]_Z8991\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(188),
    D => \GRLFPC20.FPO.FRAC\(43),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[189]_Z8992\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(189),
    D => \GRLFPC20.FPO.FRAC\(42),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[190]_Z8993\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(190),
    D => \GRLFPC20.FPO.FRAC\(41),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[191]_Z8994\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(191),
    D => \GRLFPC20.FPO.FRAC\(40),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[192]_Z8995\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(192),
    D => \GRLFPC20.FPO.FRAC\(39),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[193]_Z8996\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(193),
    D => \GRLFPC20.FPO.FRAC\(38),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[194]_Z8997\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(194),
    D => \GRLFPC20.FPO.FRAC\(37),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[195]_Z8998\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(195),
    D => \GRLFPC20.FPO.FRAC\(36),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[166]_Z8999\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(166),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(166),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[167]_Z9000\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(167),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(167),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[168]_Z9001\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(168),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(168),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[169]_Z9002\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(169),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(169),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[170]_Z9003\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(170),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(170),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[171]_Z9004\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(171),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(171),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[172]_Z9005\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(172),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(172),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[173]_Z9006\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(173),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(173),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[174]_Z9007\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(174),
    D => N_3882,
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[175]_Z9008\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(175),
    D => N_3881,
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[176]_Z9009\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(176),
    D => N_3880,
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[177]_Z9010\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(177),
    D => \GRLFPC20.FPO.FRAC\(54),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[178]_Z9011\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(178),
    D => \GRLFPC20.FPO.FRAC\(53),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[179]_Z9012\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(179),
    D => \GRLFPC20.FPO.FRAC\(52),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[180]_Z9013\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(180),
    D => \GRLFPC20.FPO.FRAC\(51),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZTREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[151]_Z9014\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(151),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(151),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[152]_Z9015\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(152),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(152),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[153]_Z9016\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(153),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(153),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[154]_Z9017\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(154),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(154),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[155]_Z9018\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(155),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(155),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[156]_Z9019\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(156),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(156),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[157]_Z9020\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(157),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(157),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[158]_Z9021\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(158),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(158),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[159]_Z9022\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(159),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(159),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[160]_Z9023\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(160),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(160),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[161]_Z9024\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(161),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(161),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[162]_Z9025\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(162),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(162),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[163]_Z9026\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(163),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(163),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[164]_Z9027\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(164),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(164),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[165]_Z9028\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(165),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(165),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[136]_Z9029\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(136),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(136),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[137]_Z9030\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(137),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(137),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[138]_Z9031\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(138),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(138),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[139]_Z9032\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(139),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(139),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[140]_Z9033\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(140),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(140),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[141]_Z9034\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(141),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(141),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[142]_Z9035\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(142),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(142),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[143]_Z9036\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(143),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(143),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[144]_Z9037\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(144),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(144),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[145]_Z9038\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(145),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(145),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[146]_Z9039\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(146),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(146),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[147]_Z9040\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(147),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(147),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[148]_Z9041\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(148),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(148),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[149]_Z9042\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(149),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(149),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[150]_Z9043\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(150),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(150),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[121]_Z9044\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(121),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(121),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[122]_Z9045\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(122),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(122),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[123]_Z9046\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(123),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(123),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[124]_Z9047\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(124),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(124),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[125]_Z9048\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(125),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(125),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[126]_Z9049\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(126),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(126),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[127]_Z9050\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(127),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(127),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[128]_Z9051\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(128),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(128),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[129]_Z9052\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(129),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(129),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[130]_Z9053\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(130),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(130),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[131]_Z9054\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(131),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(131),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[132]_Z9055\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(132),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(132),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[133]_Z9056\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(133),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(133),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[134]_Z9057\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(134),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(134),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[135]_Z9058\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(135),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(135),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[106]_Z9059\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(106),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[107]_Z9060\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(107),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[108]_Z9061\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(108),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[109]_Z9062\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(109),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[110]_Z9063\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(110),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[111]_Z9064\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(111),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[112]_Z9065\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(112),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[113]_Z9066\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(113),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[114]_Z9067\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(114),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(114),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[115]_Z9068\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(115),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(115),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[116]_Z9069\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(116),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(116),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[117]_Z9070\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(117),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(117),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[118]_Z9071\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(118),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(118),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[119]_Z9072\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(119),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(119),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[120]_Z9073\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(120),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(120),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[91]_Z9074\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(91),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[92]_Z9075\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(92),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[93]_Z9076\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(93),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[94]_Z9077\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(94),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[95]_Z9078\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(95),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[96]_Z9079\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(96),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[97]_Z9080\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(97),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[98]_Z9081\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(98),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[99]_Z9082\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(99),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[100]_Z9083\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(100),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[101]_Z9084\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(101),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[102]_Z9085\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(102),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[103]_Z9086\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(103),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[104]_Z9087\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(104),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[105]_Z9088\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(105),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[76]_Z9089\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(76),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[77]_Z9090\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(77),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[78]_Z9091\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(78),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[79]_Z9092\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(79),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[80]_Z9093\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(80),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[81]_Z9094\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(81),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[82]_Z9095\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(82),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[83]_Z9096\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(83),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[84]_Z9097\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(84),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[85]_Z9098\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(85),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[86]_Z9099\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(86),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[87]_Z9100\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(87),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[88]_Z9101\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(88),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[89]_Z9102\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(89),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[90]_Z9103\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(90),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[61]_Z9104\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(61),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[62]_Z9105\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(62),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[63]_Z9106\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(63),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[64]_Z9107\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(64),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[65]_Z9108\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(65),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[66]_Z9109\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(66),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[67]_Z9110\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(67),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[68]_Z9111\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(68),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[69]_Z9112\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(69),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[70]_Z9113\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(70),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[71]_Z9114\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(71),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[72]_Z9115\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(72),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[73]_Z9116\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(73),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[74]_Z9117\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(74),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[75]_Z9118\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(75),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[46]_Z9119\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(46),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[47]_Z9120\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(47),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[48]_Z9121\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(48),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[49]_Z9122\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(49),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[50]_Z9123\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(50),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[51]_Z9124\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(51),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[52]_Z9125\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(52),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[53]_Z9126\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(53),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[54]_Z9127\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(54),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[55]_Z9128\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(55),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[56]_Z9129\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(56),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[57]_Z9130\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(57),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[58]_Z9131\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(58),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[59]_Z9132\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(59),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[60]_Z9133\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(60),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[31]_Z9134\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(31),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[32]_Z9135\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(32),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[33]_Z9136\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(33),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[34]_Z9137\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(34),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[35]_Z9138\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(35),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[36]_Z9139\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(36),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[37]_Z9140\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(37),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[38]_Z9141\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(38),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[39]_Z9142\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(39),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[40]_Z9143\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(40),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[41]_Z9144\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(41),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[42]_Z9145\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(42),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[43]_Z9146\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(43),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[44]_Z9147\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(44),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[45]_Z9148\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(45),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[16]_Z9149\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(16),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[17]_Z9150\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(17),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[18]_Z9151\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(18),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[19]_Z9152\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(19),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[20]_Z9153\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(20),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[21]_Z9154\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(21),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[22]_Z9155\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(22),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[23]_Z9156\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(23),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[24]_Z9157\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(24),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[25]_Z9158\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(25),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[26]_Z9159\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(26),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[27]_Z9160\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(27),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[28]_Z9161\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(28),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[29]_Z9162\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(29),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[30]_Z9163\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(30),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[1]_Z9164\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(1),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[2]_Z9165\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(2),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[3]_Z9166\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(3),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[4]_Z9167\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(4),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[5]_Z9168\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(5),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[6]_Z9169\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(6),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[7]_Z9170\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(7),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[8]_Z9171\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(8),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[9]_Z9172\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(9),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[10]_Z9173\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(10),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[11]_Z9174\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(11),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[12]_Z9175\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(12),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[13]_Z9176\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(13),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[14]_Z9177\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(14),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[15]_Z9178\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(15),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[0]_Z9179\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(0),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
\GRLFPC20.RST_I\: INV port map (
    I => rst,
    O => RST_I);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CRY_0_CY_RNO\: LUT3 
generic map(
  INIT => X"B8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(35),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.MIXOIN\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_11_Z9182\: LUT2 
generic map(
  INIT => X"9"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(233),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(246),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_11\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_10_Z9183\: LUT2 
generic map(
  INIT => X"9"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(234),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(247),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_10\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_9_Z9184\: LUT2 
generic map(
  INIT => X"9"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(235),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(248),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_9\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_8_Z9185\: LUT2 
generic map(
  INIT => X"9"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(236),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(249),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_8\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_7_Z9186\: LUT2 
generic map(
  INIT => X"9"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(237),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(250),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_7\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_6_Z9187\: LUT2 
generic map(
  INIT => X"9"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(238),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(251),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_6\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_5_Z9188\: LUT2 
generic map(
  INIT => X"9"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(239),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(252),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_5\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_4_Z9189\: LUT2 
generic map(
  INIT => X"9"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(240),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(253),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_4\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_3_Z9190\: LUT2 
generic map(
  INIT => X"9"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(241),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(254),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_2_Z9191\: LUT2 
generic map(
  INIT => X"9"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(242),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(255),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_1_Z9192\: LUT2 
generic map(
  INIT => X"9"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(243),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(256),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_AXB_0\: LUT2 
generic map(
  INIT => X"9"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(257),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_I\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[235]\: LUT5 
generic map(
  INIT => X"F0AACCCC"
)
port map (
  I0 => \GRLFPC20.FPO.EXP\(9),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8581\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(248),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(235));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[236]\: LUT5 
generic map(
  INIT => X"F0AACCCC"
)
port map (
  I0 => \GRLFPC20.FPO.EXP\(8),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8580\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(249),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(236));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[234]\: LUT5 
generic map(
  INIT => X"F0AACCCC"
)
port map (
  I0 => \GRLFPC20.FPO.EXP\(10),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8582\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(247),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(234));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[235]_Z9197\: FDR port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(235),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(235),
    C => clk,
    R => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_4\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[236]_Z9198\: FDR port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(236),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(236),
    C => clk,
    R => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_4\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[234]_Z9199\: FDR port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(234),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(234),
    C => clk,
    R => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_4\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[233]_Z9200\: FDR port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(233),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(233),
    C => clk,
    R => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_4\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[232]_Z9201\: FDR port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(232),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(232),
    C => clk,
    R => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_4\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNO[71]\: LUT5 
generic map(
  INIT => X"FABAFAFA"
)
port map (
  I0 => \GRLFPC20.FPI.START\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14_2\(77),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.TEMP_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(63),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.UN38_PCTRL_NEW_I_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[257]_Z9203\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(257),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(257),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[256]_Z9204\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(256),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(256),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[255]_Z9205\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(255),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(255),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[254]_Z9206\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(254),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(254),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[253]_Z9207\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(253),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(253),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[252]_Z9208\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(252),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(252),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[251]_Z9209\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(251),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(251),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[250]_Z9210\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(250),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(250),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[245]_Z9211\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(245),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(245),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH[246]_Z9212\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(246),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(246),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[40]_Z9213\: FDE port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(40),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_21\(40),
    C => clk,
    CE => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_21_0[40]\: LUT2 
generic map(
  INIT => X"E"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1776\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_21_0_1_TZ\(40),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_21\(40));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH[254]_Z9215\: LUT3 
generic map(
  INIT => X"E4"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8781\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41\(254),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(254));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_0[257]\: LUT5 
generic map(
  INIT => X"F0CCAAAA"
)
port map (
  I0 => \GRLFPC20.FPO.EXP\(0),
  I1 => \GRLFPC20.FPO.EXP\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_1[257]\: LUT5 
generic map(
  INIT => X"FCAC5C0C"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  I1 => \GRLFPC20.FPI.OP1\(52),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => rfo1_data1(23),
  I4 => rfo2_data1(23),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[257]\: MUXF7 port map (
    I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0\,
    I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1\,
    S => \GRLFPC20.FPI.LDOP\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(257));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_0[256]\: LUT5 
generic map(
  INIT => X"F0CCAAAA"
)
port map (
  I0 => \GRLFPC20.FPO.EXP\(1),
  I1 => \GRLFPC20.FPO.EXP\(2),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(243),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_1[256]\: LUT5 
generic map(
  INIT => X"FCAC5C0C"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  I1 => \GRLFPC20.FPI.OP1\(53),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => rfo1_data1(24),
  I4 => rfo2_data1(24),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[256]\: MUXF7 port map (
    I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_0\,
    I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_0\,
    S => \GRLFPC20.FPI.LDOP\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(256));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_0[255]\: LUT5 
generic map(
  INIT => X"F0CCAAAA"
)
port map (
  I0 => \GRLFPC20.FPO.EXP\(2),
  I1 => \GRLFPC20.FPO.EXP\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(242),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_1[255]\: LUT5 
generic map(
  INIT => X"FCAC5C0C"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  I1 => \GRLFPC20.FPI.OP1\(54),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => rfo1_data1(25),
  I4 => rfo2_data1(25),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[255]\: MUXF7 port map (
    I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_1\,
    I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_1\,
    S => \GRLFPC20.FPI.LDOP\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(255));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_0[252]\: LUT5 
generic map(
  INIT => X"F0CCAAAA"
)
port map (
  I0 => \GRLFPC20.FPO.EXP\(5),
  I1 => \GRLFPC20.FPO.EXP\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(239),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_1[252]\: LUT5 
generic map(
  INIT => X"CFCAC5C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  I1 => \GRLFPC20.FPI.OP1\(60),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => rfo1_data1(25),
  I4 => rfo2_data1(25),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[252]\: MUXF7 port map (
    I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_2\,
    I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_2\,
    S => \GRLFPC20.FPI.LDOP\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(252));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_0[251]\: LUT5 
generic map(
  INIT => X"F0CCAAAA"
)
port map (
  I0 => \GRLFPC20.FPO.EXP\(6),
  I1 => \GRLFPC20.FPO.EXP\(7),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(238),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_1[251]\: LUT5 
generic map(
  INIT => X"CFCAC5C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  I1 => \GRLFPC20.FPI.OP1\(61),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => rfo1_data1(26),
  I4 => rfo2_data1(26),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[251]\: MUXF7 port map (
    I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_3\,
    I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_3\,
    S => \GRLFPC20.FPI.LDOP\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(251));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_0[250]\: LUT5 
generic map(
  INIT => X"F0CCAAAA"
)
port map (
  I0 => \GRLFPC20.FPO.EXP\(7),
  I1 => \GRLFPC20.FPO.EXP\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(237),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_4\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_1[250]\: LUT5 
generic map(
  INIT => X"CFCAC5C0"
)
port map (
  I0 => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
  I1 => \GRLFPC20.FPI.OP1\(62),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  I3 => rfo1_data1(27),
  I4 => rfo2_data1(27),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_4\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[250]\: MUXF7 port map (
    I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_4\,
    I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_4\,
    S => \GRLFPC20.FPI.LDOP\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(250));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[245]\: LUT5 
generic map(
  INIT => X"30222222"
)
port map (
  I0 => N_3812,
  I1 => \GRLFPC20.FPI.LDOP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(232),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(245));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[246]\: LUT6 
generic map(
  INIT => X"0F000C0C0A0A0A0A"
)
port map (
  I0 => N_3811,
  I1 => N_3812,
  I2 => \GRLFPC20.FPI.LDOP\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(233),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(246));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[232]\: LUT6 
generic map(
  INIT => X"FF00AAAA30303030"
)
port map (
  I0 => N_3812,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(232),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(245),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(232));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[233]\: LUT6 
generic map(
  INIT => X"FF00AAAA30303030"
)
port map (
  I0 => N_3811,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(233),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(246),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(233));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_RNO_0[19]\: LUT6 
generic map(
  INIT => X"CCCC00A000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9637_I\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9666_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3I0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_RNO_1[19]\: LUT6 
generic map(
  INIT => X"AAAA00C000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9666_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3I1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_8_RNO[19]\: MUXF7 port map (
    I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3I0\,
    I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3I1\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_3\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_RNO_0[33]\: LUT6 
generic map(
  INIT => X"DC00CC00CC00CC00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_52\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9919_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1I0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_RNO_1[33]\: LUT6 
generic map(
  INIT => X"0000000088000800"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1I1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_6_RNO[33]\: MUXF7 port map (
    I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1I0\,
    I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1I1\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(33));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_RNO_0[52]\: LUT6 
generic map(
  INIT => X"2000000000000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_717\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10025_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1I0_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_RNO_1[52]\: LUT6 
generic map(
  INIT => X"0044004400030300"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_715\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1I1_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_11_RNO[52]\: MUXF7 port map (
    I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1I0_0\,
    I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1I1_0\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_RNO_0[53]\: LUT6 
generic map(
  INIT => X"EEEAAAAAEAAAAAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7\(53),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A22_11_0\(53),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9I0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_RNO_1[53]\: LUT6 
generic map(
  INIT => X"FCF0F0FAFCF0F0F0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10284\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10694_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_7\(53),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9I1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_RNO[53]\: MUXF7 port map (
    I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9I0\,
    I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9I1\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_9\(53));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_0[239]\: LUT5 
generic map(
  INIT => X"CFC0AFA0"
)
port map (
  I0 => \GRLFPC20.FPI.OP2\(57),
  I1 => \GRLFPC20.FPI.OP2\(60),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(239),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_5\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_1[239]\: LUT5 
generic map(
  INIT => X"F0CCAACC"
)
port map (
  I0 => \GRLFPC20.FPO.EXP\(5),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(252),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(27),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_5\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[239]\: MUXF7 port map (
    I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_5\,
    I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_5\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_3\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(239));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_0[240]\: LUT5 
generic map(
  INIT => X"CFC0AFA0"
)
port map (
  I0 => \GRLFPC20.FPI.OP2\(56),
  I1 => \GRLFPC20.FPI.OP2\(59),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(240),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_6\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_1[240]\: LUT5 
generic map(
  INIT => X"F0CCAACC"
)
port map (
  I0 => \GRLFPC20.FPO.EXP\(4),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(253),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(27),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_6\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[240]\: MUXF7 port map (
    I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_6\,
    I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_6\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_3\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(240));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_0[242]\: LUT5 
generic map(
  INIT => X"CFC0AFA0"
)
port map (
  I0 => \GRLFPC20.FPI.OP2\(54),
  I1 => \GRLFPC20.FPI.OP2\(57),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(242),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_7\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_1[242]\: LUT5 
generic map(
  INIT => X"F0CCAACC"
)
port map (
  I0 => \GRLFPC20.FPO.EXP\(2),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(255),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(27),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_7\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[242]\: MUXF7 port map (
    I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_7\,
    I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_7\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_3\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(242));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_0[56]\: LUT6 
generic map(
  INIT => X"3333F0F055005500"
)
port map (
  I0 => \GRLFPC20.FPI.LDOP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8691\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(114),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(172),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_1[56]\: LUT5 
generic map(
  INIT => X"0A0CFA0C"
)
port map (
  I0 => N_3825,
  I1 => N_3826,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_25\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[56]\: MUXF7 port map (
    I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I0\,
    I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I1\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(56));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_0[243]\: LUT5 
generic map(
  INIT => X"CFC0AFA0"
)
port map (
  I0 => \GRLFPC20.FPI.OP2\(53),
  I1 => \GRLFPC20.FPI.OP2\(56),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(243),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_8\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_1[243]\: LUT5 
generic map(
  INIT => X"F0CCAACC"
)
port map (
  I0 => \GRLFPC20.FPO.EXP\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(256),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(27),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_8\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[243]\: MUXF7 port map (
    I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_8\,
    I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_8\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_3\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(243));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_0[238]\: LUT5 
generic map(
  INIT => X"CFC0AFA0"
)
port map (
  I0 => \GRLFPC20.FPI.OP2\(58),
  I1 => \GRLFPC20.FPI.OP2\(61),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(238),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_9\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_1[238]\: LUT5 
generic map(
  INIT => X"F0CCAACC"
)
port map (
  I0 => \GRLFPC20.FPO.EXP\(6),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(251),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(27),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_9\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[238]\: MUXF7 port map (
    I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_9\,
    I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_9\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_3\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(238));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_0[241]\: LUT5 
generic map(
  INIT => X"CFC0AFA0"
)
port map (
  I0 => \GRLFPC20.FPI.OP2\(55),
  I1 => \GRLFPC20.FPI.OP2\(58),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(241),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_10\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_1[241]\: LUT5 
generic map(
  INIT => X"F0CCAACC"
)
port map (
  I0 => \GRLFPC20.FPO.EXP\(3),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(254),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(27),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_10\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[241]\: MUXF7 port map (
    I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_10\,
    I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_10\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_3\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(241));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_0[237]\: LUT5 
generic map(
  INIT => X"CFC0AFA0"
)
port map (
  I0 => \GRLFPC20.FPI.OP2\(59),
  I1 => \GRLFPC20.FPI.OP2\(62),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(237),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_11\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_1[237]\: LUT5 
generic map(
  INIT => X"F0CCAACC"
)
port map (
  I0 => \GRLFPC20.FPO.EXP\(7),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(250),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(27),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_11\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[237]\: MUXF7 port map (
    I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI0_11\,
    I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATHI1_11\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_N_3\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(237));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_0[38]\: LUT5 
generic map(
  INIT => X"33F0AAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7879\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8709\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I0_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_1[38]\: LUT6 
generic map(
  INIT => X"F0F0AAAAFF00CCCC"
)
port map (
  I0 => \GRLFPC20.FPO.FRAC\(18),
  I1 => \GRLFPC20.FPO.FRAC\(19),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(38),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I1_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[38]\: MUXF7 port map (
    I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I0_0\,
    I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I1_0\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(38));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_0[35]\: LUT5 
generic map(
  INIT => X"33F0AAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7882\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8712\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I0_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_1[35]\: LUT6 
generic map(
  INIT => X"F0F0AAAAFF00CCCC"
)
port map (
  I0 => \GRLFPC20.FPO.FRAC\(21),
  I1 => \GRLFPC20.FPO.FRAC\(22),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(35),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I1_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[35]\: MUXF7 port map (
    I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I0_1\,
    I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I1_1\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(35));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_0[34]\: LUT5 
generic map(
  INIT => X"33F0AAAA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7883\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8713\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_7_MUX\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I0_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO_1[34]\: LUT6 
generic map(
  INIT => X"F0F0AAAAFF00CCCC"
)
port map (
  I0 => \GRLFPC20.FPO.FRAC\(22),
  I1 => \GRLFPC20.FPO.FRAC\(23),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(34),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I1_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNO[34]\: MUXF7 port map (
    I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I0_2\,
    I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1I1_2\,
    S => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH1\(34));
\GRLFPC20.R.A.RF1REN_RNO[1]\: LUT5 
generic map(
  INIT => X"0202FF00"
)
port map (
  I0 => \GRLFPC20.COMB.RS1V_1\,
  I1 => \GRLFPC20.COMB.V.A.RF1REN_1_115_I_0\,
  I2 => \GRLFPC20.COMB.LOCKGEN.LOCKI\,
  I3 => \GRLFPC20.R.A.RF1REN\(1),
  I4 => holdn,
  O => \GRLFPC20.N_2994_I_0\);
\GRLFPC20.COMB.V.A.RF1REN_1[2]\: LUT6 
generic map(
  INIT => X"00C400C4FFFF0000"
)
port map (
  I0 => cpi_d_inst(0),
  I1 => \GRLFPC20.N_1583\,
  I2 => \GRLFPC20.COMB.RS2D_1\,
  I3 => \GRLFPC20.COMB.LOCKGEN.LOCKI\,
  I4 => \GRLFPC20.R.A.RF1REN\(2),
  I5 => holdn,
  O => \GRLFPC20.COMB.V.A.RF1REN_1_0\(2));
\GRLFPC20.COMB.RS1_1_0_0[1]_Z9285\: LUT6 
generic map(
  INIT => X"ACA0ACA0FFFF0000"
)
port map (
  I0 => cpi_d_inst(15),
  I1 => cpi_d_inst(26),
  I2 => \GRLFPC20.N_1583\,
  I3 => \GRLFPC20.RS1V_0_SQMUXA\,
  I4 => \GRLFPC20.R.A.RS1\(1),
  I5 => holdn,
  O => \GRLFPC20.COMB.RS1_1_0_0\(1));
\GRLFPC20.COMB.RS1_1_0_0[2]_Z9286\: LUT6 
generic map(
  INIT => X"ACA0ACA0FFFF0000"
)
port map (
  I0 => cpi_d_inst(16),
  I1 => cpi_d_inst(27),
  I2 => \GRLFPC20.N_1583\,
  I3 => \GRLFPC20.RS1V_0_SQMUXA\,
  I4 => \GRLFPC20.R.A.RS1\(2),
  I5 => holdn,
  O => \GRLFPC20.COMB.RS1_1_0_0\(2));
\GRLFPC20.COMB.RS1_1_0_0[3]_Z9287\: LUT6 
generic map(
  INIT => X"ACA0ACA0FFFF0000"
)
port map (
  I0 => cpi_d_inst(17),
  I1 => cpi_d_inst(28),
  I2 => \GRLFPC20.N_1583\,
  I3 => \GRLFPC20.RS1V_0_SQMUXA\,
  I4 => \GRLFPC20.R.A.RS1\(3),
  I5 => holdn,
  O => \GRLFPC20.COMB.RS1_1_0_0\(3));
\GRLFPC20.COMB.RS1_1_0_0[4]_Z9288\: LUT6 
generic map(
  INIT => X"ACA0ACA0FFFF0000"
)
port map (
  I0 => cpi_d_inst(18),
  I1 => cpi_d_inst(29),
  I2 => \GRLFPC20.N_1583\,
  I3 => \GRLFPC20.RS1V_0_SQMUXA\,
  I4 => \GRLFPC20.R.A.RS1\(4),
  I5 => holdn,
  O => \GRLFPC20.COMB.RS1_1_0_0\(4));
\GRLFPC20.COMB.RS2_1[2]\: LUT4 
generic map(
  INIT => X"88F0"
)
port map (
  I0 => cpi_d_inst(2),
  I1 => \GRLFPC20.N_1583\,
  I2 => \GRLFPC20.R.A.RS2\(2),
  I3 => holdn,
  O => \GRLFPC20.COMB.RS2_1_0\(2));
\GRLFPC20.COMB.RS2_1[1]\: LUT4 
generic map(
  INIT => X"88F0"
)
port map (
  I0 => cpi_d_inst(1),
  I1 => \GRLFPC20.N_1583\,
  I2 => \GRLFPC20.R.A.RS2\(1),
  I3 => holdn,
  O => \GRLFPC20.COMB.RS2_1_0\(1));
\GRLFPC20.COMB.RS2_1[3]\: LUT4 
generic map(
  INIT => X"88F0"
)
port map (
  I0 => cpi_d_inst(3),
  I1 => \GRLFPC20.N_1583\,
  I2 => \GRLFPC20.R.A.RS2\(3),
  I3 => holdn,
  O => \GRLFPC20.COMB.RS2_1_0\(3));
\GRLFPC20.COMB.RS2_1[4]\: LUT4 
generic map(
  INIT => X"88F0"
)
port map (
  I0 => cpi_d_inst(4),
  I1 => \GRLFPC20.N_1583\,
  I2 => \GRLFPC20.R.A.RS2\(4),
  I3 => holdn,
  O => \GRLFPC20.COMB.RS2_1_0\(4));
\GRLFPC20.COMB.RS2_1DUP[0]_Z9293\: LUT4 
generic map(
  INIT => X"88F0"
)
port map (
  I0 => cpi_d_inst(0),
  I1 => \GRLFPC20.N_1583\,
  I2 => \GRLFPC20.R.A.RS2\(0),
  I3 => holdn,
  O => \GRLFPC20.COMB.RS2_1DUP\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_RNO[8]\: LUT6 
generic map(
  INIT => X"FDFCFDFCFFFF0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(2),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(21),
  I3 => \GRLFPC20.R.FSR.RD\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(8),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.TEMP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.U_RDN_1_5599\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_RNO[9]\: LUT5 
generic map(
  INIT => X"FEFEFF00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(21),
  I2 => \GRLFPC20.R.FSR.RD\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(9),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.TEMP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_11210_I_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_RNI214P1[13]\: LUT6 
generic map(
  INIT => X"44044404FFFF0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(38),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(39),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(13),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(40),
  I4 => \GRLFPC20.R.I.CC\(1),
  I5 => \GRLFPC20.N_2102\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_587_I_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_RNI104P1[13]\: LUT6 
generic map(
  INIT => X"44404440FFFF0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(38),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(39),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(13),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(40),
  I4 => \GRLFPC20.R.I.CC\(0),
  I5 => \GRLFPC20.N_2102\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_589_I_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNO[65]\: LUT6 
generic map(
  INIT => X"FFFFFFFFE0F0FFFF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.ENTRYPOINT\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(66),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(67),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(68),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(64),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_2_0_E\(65));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNO[69]\: LUT6 
generic map(
  INIT => X"FFFFFFFF1F0F1000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.ENTRYPOINT\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(66),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(67),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(69),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(64),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_E_0_E\(69));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNO[73]\: LUT4 
generic map(
  INIT => X"0073"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.ENTRYPOINT\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(66),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(67),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN3_NOTRESETORUNIMP_0_E\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNO[77]\: LUT6 
generic map(
  INIT => X"000000004CCC0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.OPREXCSHFT.UN3_OPREXC\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14_2\(77),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1\(5),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(46),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14_0_E\(77));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_RNO[6]\: LUT5 
generic map(
  INIT => X"00002070"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.U_RDN_1\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_10\(10),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(8),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(9),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_16_0_E\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_RNO[5]\: LUT4 
generic map(
  INIT => X"0027"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.TEMP\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.U_RDN_1\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(8),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(9),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.UN53_SCTRL_NEW_I_0_E\);
\GRLFPC20.R.MK.HOLDN1_RNO\: LUT2 
generic map(
  INIT => X"D"
)
port map (
  I0 => \GRLFPC20.R.MK.RST2\,
  I1 => RST_I,
  O => \GRLFPC20.R.MK.RST2_I_E\);
\GRLFPC20.R.A.RS2[0]_Z9305\: FD port map (
    Q => \GRLFPC20.R.A.RS2\(0),
    D => \GRLFPC20.COMB.RS2_1DUP\(0),
    C => clk);
\GRLFPC20.R.A.RS2[4]_Z9306\: FD port map (
    Q => \GRLFPC20.R.A.RS2\(4),
    D => \GRLFPC20.COMB.RS2_1_0\(4),
    C => clk);
\GRLFPC20.R.A.RS2[3]_Z9307\: FD port map (
    Q => \GRLFPC20.R.A.RS2\(3),
    D => \GRLFPC20.COMB.RS2_1_0\(3),
    C => clk);
\GRLFPC20.R.A.RS2[1]_Z9308\: FD port map (
    Q => \GRLFPC20.R.A.RS2\(1),
    D => \GRLFPC20.COMB.RS2_1_0\(1),
    C => clk);
\GRLFPC20.R.A.RS2[2]_Z9309\: FD port map (
    Q => \GRLFPC20.R.A.RS2\(2),
    D => \GRLFPC20.COMB.RS2_1_0\(2),
    C => clk);
\GRLFPC20.R.A.RS1[4]_Z9310\: FD port map (
    Q => \GRLFPC20.R.A.RS1\(4),
    D => \GRLFPC20.COMB.RS1_1_0_0\(4),
    C => clk);
\GRLFPC20.R.A.RS1[3]_Z9311\: FD port map (
    Q => \GRLFPC20.R.A.RS1\(3),
    D => \GRLFPC20.COMB.RS1_1_0_0\(3),
    C => clk);
\GRLFPC20.R.A.RS1[2]_Z9312\: FD port map (
    Q => \GRLFPC20.R.A.RS1\(2),
    D => \GRLFPC20.COMB.RS1_1_0_0\(2),
    C => clk);
\GRLFPC20.R.A.RS1[1]_Z9313\: FD port map (
    Q => \GRLFPC20.R.A.RS1\(1),
    D => \GRLFPC20.COMB.RS1_1_0_0\(1),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[65]_Z9314\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_2_0_E\(65),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[68]_Z9315\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(68),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN2_NOTDECODEDUNIMP_0_E\,
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[69]_Z9316\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(69),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_E_0_E\(69),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL[1]_Z9317\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(1),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_5_0_E\(1),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL[2]_Z9318\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(2),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_4_0_E\(2),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL[0]_Z9319\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(0),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_6_0_E\(0),
    C => clk);
\GRLFPC20.R.MK.LDOP_Z9320\: FD port map (
    Q => \GRLFPC20.R.MK.LDOP\,
    D => \GRLFPC20.RIN.MK.LDOP_0_E\,
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[77]_Z9321\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(77),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14_0_E\(77),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL[73]_Z9322\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(73),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN3_NOTRESETORUNIMP_0_E\,
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL[6]_Z9323\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(6),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_16_0_E\(6),
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL[5]_Z9324\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(5),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.UN53_SCTRL_NEW_I_0_E\,
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL[9]_Z9325\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(9),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_11210_I_0\,
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL[8]_Z9326\: FD port map (
    Q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(8),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.U_RDN_1_5599\,
    C => clk);
\GRLFPC20.R.A.RF1REN[2]_Z9327\: FD port map (
    Q => \GRLFPC20.R.A.RF1REN\(2),
    D => \GRLFPC20.COMB.V.A.RF1REN_1_0\(2),
    C => clk);
\GRLFPC20.R.A.RF1REN[1]_Z9328\: FD port map (
    Q => \GRLFPC20.R.A.RF1REN\(1),
    D => \GRLFPC20.N_2994_I_0\,
    C => clk);
\GRLFPC20.R.I.CC[0]_Z9329\: FD port map (
    Q => \GRLFPC20.R.I.CC\(0),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_589_I_0\,
    C => clk);
\GRLFPC20.R.I.CC[1]_Z9330\: FD port map (
    Q => \GRLFPC20.R.I.CC\(1),
    D => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_587_I_0\,
    C => clk);
\GRLFPC20.R.MK.HOLDN1_Z9331\: FD port map (
    Q => \GRLFPC20.R.MK.HOLDN1\,
    D => \GRLFPC20.R.MK.RST2_I_E\,
    C => clk);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_23_LUT6_2[52]\: LUT6_2 
generic map(
  INIT => X"0000000000200000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_765\,
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2129\,
  O5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2772\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_3_LUT6_2[3]\: LUT6_2 
generic map(
  INIT => X"0000000010000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2563\,
  O5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10243_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_14_LUT6_2[57]\: LUT6_2 
generic map(
  INIT => X"0000000000000080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1019_1\,
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10619\,
  O5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A24_0\(59));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_13_LUT6_2[36]\: LUT6_2 
generic map(
  INIT => X"0000000000000010"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10035\,
  O5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2774\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_3_2_LUT6_2[19]\: LUT6_2 
generic map(
  INIT => X"0000010100001100"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_3_2\(19),
  O5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2601\);
\GRLFPC20.COMB.V.I.EXEC_5_IV_LUT6_2\: LUT6_2 
generic map(
  INIT => X"FFFEFFFF01000100"
)
port map (
  I0 => cpi_flush,
  I1 => cpi_x_annul,
  I2 => cpi_x_trap,
  I3 => \GRLFPC20.R.X.FPOP\,
  I4 => \GRLFPC20.R.X.SEQERR\,
  I5 => \GRLFPC20.R.I.EXEC\,
  O6 => \GRLFPC20.COMB.V.I.EXEC_5\,
  O5 => \GRLFPC20.V.I.EXEC_0_SQMUXA\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_0_A2_LUT6_2[46]\: LUT6_2 
generic map(
  INIT => X"0000000000001200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2206\,
  O5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9971\);
\GRLFPC20.COMB.UN1_V.STATE_LUT6_2\: LUT6_2 
generic map(
  INIT => X"0000000000050003"
)
port map (
  I0 => \GRLFPC20.R.STATE\(0),
  I1 => \GRLFPC20.R.X.SEQERR\,
  I2 => \GRLFPC20.N_2000\,
  I3 => \GRLFPC20.N_2015\,
  I4 => \GRLFPC20.V.STATE_2_SQMUXA\,
  I5 => \GRLFPC20.COMB.V.STATE_9\(1),
  O6 => \GRLFPC20.N_2074\,
  O5 => \GRLFPC20.COMB.V.STATE_9_I\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14_2_LUT6_2_RNIU2NI1[77]\: LUT6_2 
generic map(
  INIT => X"FFFDFFFFFFFDFFFD"
)
port map (
  I0 => rst,
  I1 => \GRLFPC20.R.MK.LDOP\,
  I2 => \GRLFPC20.R.MK.RST\,
  I3 => \GRLFPC20.R.MK.RST2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14\(77),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14_2\(77),
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB_I\,
  O5 => \GRLFPC20.FPI.LDOP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_I_A2_4_LUT6_2[0]\: LUT6_2 
generic map(
  INIT => X"0000000100010001"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXCEP_1_I_A2_4\(0),
  O5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_2_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12.Z_AXB1_LUT6_2\: LUT6_2 
generic map(
  INIT => X"A5C3FFFF5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.SI_12\(45),
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12.Z_AXB1\,
  O5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8.Z_AXB2_LUT6_2\: LUT6_2 
generic map(
  INIT => X"C3A5FFFF3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.SI_65\(48),
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8.Z_AXB2\,
  O5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18.Z_AXB1_LUT6_2\: LUT6_2 
generic map(
  INIT => X"C3A5FFFF3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.SI_18\(39),
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18.Z_AXB1\,
  O5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21.Z_AXB2_LUT6_2\: LUT6_2 
generic map(
  INIT => X"A5C3FFFF5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.SI_78\(35),
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21.Z_AXB2\,
  O5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_AXB1_LUT6_2\: LUT6_2 
generic map(
  INIT => X"33A5FFFFCC5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.UN255_TEMP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.SI_30\(27),
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_AXB1\,
  O5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_AXB1_LUT6_2\: LUT6_2 
generic map(
  INIT => X"A5C3FFFF5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.SI_32\(25),
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_AXB1\,
  O5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.CIN_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_AXB1_LUT6_2\: LUT6_2 
generic map(
  INIT => X"C3A5FFFF3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.SI_34\(23),
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_AXB1\,
  O5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.CIN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36.Z_AXB2_LUT6_2\: LUT6_2 
generic map(
  INIT => X"C3A5FFFF3C5A0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.SI_93\(20),
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36.Z_AXB2\,
  O5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45.Z_AXB1_LUT6_2\: LUT6_2 
generic map(
  INIT => X"A5C3FFFF5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.SI_45\(12),
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45.Z_AXB1\,
  O5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_541_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43.Z_AXB1_LUT6_2\: LUT6_2 
generic map(
  INIT => X"A5C3FFFF5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.SI_43\(14),
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43.Z_AXB1\,
  O5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_548_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39.Z_AC0_2_LUT6_2\: LUT6_2 
generic map(
  INIT => X"000000005A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.SI_39\(18),
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39.Z_AC0_2\,
  O5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_559_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48.Z_AXB0_LUT6_2\: LUT6_2 
generic map(
  INIT => X"A5C3FFFF5A3C0000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(13),
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48.Z_AXB0\,
  O5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.CIN_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_LUT6_2[4]\: LUT6_2 
generic map(
  INIT => X"0F0F555500FF3333"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8362\,
  O5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(53));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_LUT6_2[6]\: LUT6_2 
generic map(
  INIT => X"0F0F555500FF3333"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8360\,
  O5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(51));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26_LUT6_2[52]\: LUT6_2 
generic map(
  INIT => X"000000F000CC00AA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(52),
  O5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8314_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26_LUT6_2[53]\: LUT6_2 
generic map(
  INIT => X"000000AA00F000CC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  I5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  O6 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(53),
  O5 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8313_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26_LUT6_2_RNI2MC3[53]\: INV port map (
    I => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8313_I\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8313\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26_LUT6_2_RNI1LC3[52]\: INV port map (
    I => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8314_I\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8314\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_V_I_O5_INV[1]\: INV port map (
    I => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_559_I\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_559\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_V_I_O5_INV[1]\: INV port map (
    I => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_548_I\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_548\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_V_I_O5_INV[1]\: INV port map (
    I => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_541_I\,
    O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_541\);
\GRLFPC20.COMB.UN1_V.STATE_LUT6_2_RNIG4OE\: INV port map (
    I => \GRLFPC20.COMB.V.STATE_9_I\(0),
    O => \GRLFPC20.COMB.V.STATE_9\(0));
II_GND: GND port map (
    G => NN_2);
II_VCC: VCC port map (
    P => NN_3);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_LUT6_2_O6[28]\: LUT3 
generic map(
  INIT => X"1B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(28),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(29),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8659\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_LUT6_2_O5[28]\: LUT3 
generic map(
  INIT => X"27"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(28),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(27),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8660\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_LUT6_2_O6[23]\: LUT3 
generic map(
  INIT => X"1B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(23),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(24),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8664\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_LUT6_2_O5[23]\: LUT3 
generic map(
  INIT => X"1B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(14),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(15),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8673\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_LUT6_2_O6[20]\: LUT3 
generic map(
  INIT => X"1B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(20),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(21),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8667\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_LUT6_2_O5[20]\: LUT3 
generic map(
  INIT => X"27"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(20),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(19),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8668\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_LUT6_2_O6[18]\: LUT3 
generic map(
  INIT => X"1B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(18),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(19),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8669\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_LUT6_2_O5[18]\: LUT3 
generic map(
  INIT => X"27"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(18),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8670\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_LUT6_2_O6[25]\: LUT3 
generic map(
  INIT => X"1B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(25),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(26),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8662\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_LUT6_2_O5[25]\: LUT3 
generic map(
  INIT => X"27"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(25),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(24),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8663\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_LUT6_2_O6[33]\: LUT3 
generic map(
  INIT => X"1B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(33),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8654\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_LUT6_2_O5[33]\: LUT3 
generic map(
  INIT => X"27"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(53),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(52),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8635\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_LUT6_2_O6[29]\: LUT3 
generic map(
  INIT => X"27"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(30),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(29),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8658\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_LUT6_2_O5[29]\: LUT3 
generic map(
  INIT => X"1B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(30),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(31),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8657\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_LUT6_2_O6[21]\: LUT3 
generic map(
  INIT => X"1B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(21),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(22),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8666\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_LUT6_2_O5[21]\: LUT3 
generic map(
  INIT => X"1B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(22),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(23),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8665\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_LUT6_2_O6[16]\: LUT3 
generic map(
  INIT => X"1B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(16),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8671\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_LUT6_2_O5[16]\: LUT3 
generic map(
  INIT => X"1B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(15),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(16),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8672\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26_LUT6_2_O6[39]\: LUT3 
generic map(
  INIT => X"27"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8325\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8327\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(39));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26_LUT6_2_O5[39]\: LUT3 
generic map(
  INIT => X"1B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8331\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8329\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(35));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_LUT6_2_O6[47]\: LUT5 
generic map(
  INIT => X"FF330F55"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8319\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_LUT6_2_O5[47]\: LUT4 
generic map(
  INIT => X"F3F5"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8315\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_LUT6_2_O6[49]\: LUT5 
generic map(
  INIT => X"FF330F55"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8317\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_LUT6_2_O5[49]\: LUT2 
generic map(
  INIT => X"1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_S0\(3));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_LUT6_2_O6[46]\: LUT5 
generic map(
  INIT => X"FF330F55"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8320\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_LUT6_2_O5[46]\: LUT4 
generic map(
  INIT => X"F3F5"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8316\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4.Z_AXBXC3_LUT6_2_O6\: LUT3 
generic map(
  INIT => X"96"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4.Z_C3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.SI_118\(51),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4.Z_AXBXC3_LUT6_2_O5\: LUT3 
generic map(
  INIT => X"E8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4.Z_C3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.SI_118\(51),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(61));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_C4_LUT6_2_O6\: LUT3 
generic map(
  INIT => X"E8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_C3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.SI_134\(35),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(77));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_C4_LUT6_2_O5\: LUT3 
generic map(
  INIT => X"96"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_C3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.SI_134\(35),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(20));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19.Z_C4_LUT6_2_O6\: LUT3 
generic map(
  INIT => X"E8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.SI_133\(36),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(76));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19.Z_C4_LUT6_2_O5\: LUT3 
generic map(
  INIT => X"96"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.SI_133\(36),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18.Z_C4_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"B2E8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_C2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18.Z_C3\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_AXB2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(75));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18.Z_C4_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"6996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_C2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18.Z_C3\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17.Z_AXB2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(18));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_AXBXC3_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"96696996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14.Z_C2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.SI_71\(42),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(15));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_AXBXC3_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"EBBE8228"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14.Z_C2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.SI_71\(42),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(72));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8.Z_AXBXC3_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"6996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7.Z_C2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7.Z_AXB2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(8));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8.Z_AXBXC3_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"BE28"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7.Z_C2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7.Z_AXB2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(65));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31.Z_C4_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"EBBE8228"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_C2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.SI_87\(26),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(88));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31.Z_C4_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"96696996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_C2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.SI_87\(26),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(31));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_C4_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"EBBE8228"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.SI_85\(28),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(86));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_C4_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"96696996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.SI_85\(28),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(29));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26.Z_C4_LUT6_2_O6\: LUT3 
generic map(
  INIT => X"E8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26.Z_C3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.SI_140\(29),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(83));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26.Z_C4_LUT6_2_O5\: LUT3 
generic map(
  INIT => X"96"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26.Z_C3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.SI_140\(29),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(26));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_C4_LUT6_2_O6\: LUT3 
generic map(
  INIT => X"E8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.SI_139\(30),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(82));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_C4_LUT6_2_O5\: LUT3 
generic map(
  INIT => X"96"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.SI_139\(30),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(25));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_C4_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"EBBE8228"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22.Z_C2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.SI_79\(34),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(80));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_C4_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"96696996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22.Z_C2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.SI_79\(34),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(23));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44.Z_C4_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"EBBE8228"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.SI_100\(13),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(101));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44.Z_C4_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"96696996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.SI_100\(13),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(44));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39.Z_C4_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"EBBE8228"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.SI_95\(18),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(96));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39.Z_C4_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"96696996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.SI_95\(18),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(39));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38.Z_C4_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"FEEAA880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.SI_95\(18),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.SI_152\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(95));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38.Z_C4_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"A995566A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.SI_95\(18),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.SI_152\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(38));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50.Z_C4_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"BE28"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49.Z_AXB2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49.Z_C2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(107));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50.Z_C4_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"6996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49.Z_AXB2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49.Z_C2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(50));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49.Z_C4_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"FEEAA880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.SI_106\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.SI_163\(6),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(106));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49.Z_C4_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"A995566A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.SI_106\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.SI_163\(6),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(49));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47.Z_C4_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"BE28"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_C2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_AXB2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(104));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47.Z_C4_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"6996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_C2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_AXB2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47.Z_C3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_C4_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"FEEAA880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.SI_103\(10),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.SI_160\(9),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(103));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_C4_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"A995566A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.SI_103\(10),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.SI_160\(9),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(46));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55.Z_C4_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"FEEAA880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.SI_112\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(112));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55.Z_C4_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"A995566A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.SI_112\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55.Z_C2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8\(55));
\GRLFPC20.COMB.V.A.SEQERR_1_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"0000AACA"
)
port map (
  I0 => \GRLFPC20.COMB.V.A.AFQ_1_1\,
  I1 => \GRLFPC20.N_1138\,
  I2 => \GRLFPC20.R.STATE\(1),
  I3 => \GRLFPC20.R.STATE\(0),
  I4 => \GRLFPC20.N_1317\,
  O => \GRLFPC20.COMB.V.A.SEQERR_1\);
\GRLFPC20.COMB.V.A.SEQERR_1_LUT6_2_O5\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => \GRLFPC20.R.STATE\(1),
  I1 => \GRLFPC20.R.STATE\(0),
  O => CPO_EXC_1);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_C3_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"EDDE8448"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.SI_19\(38),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19.Z_C1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_C3_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"6996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.SI_19\(38),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19.Z_C1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20.Z_AXB2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_C3_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"FEECC880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.SI_15\(42),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_C1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.SI_72\(41),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_C3_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"C993366C"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.SI_15\(42),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_C1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.SI_72\(41),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.SI_130\(39));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12.Z_C3_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"EDDE8448"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.SI_11\(46),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12.Z_C3_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"96696996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.SI_11\(46),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.SI_127\(42));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11.Z_C3_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"FEECC880"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.SI_11\(46),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.SI_68\(45),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11.Z_C3_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"C993366C"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.SI_11\(46),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.SI_68\(45),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.SI_126\(43));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9.Z_C3_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"EBBE8228"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.SI_8\(49),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9.Z_C3_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"96696996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.SI_8\(49),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.SI_124\(45));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_C3_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"EBBE8228"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.SI_33\(24),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_C3_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"96696996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.CIN_3\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.CIN_2\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.SI_33\(24),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.SI_149\(20));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45.Z_C3_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"BEEB2882"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_544\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.SI_44\(13),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45.Z_C3_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"69969669"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_544\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.SI_44\(13),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.SI_160\(9));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37.Z_C3_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"EBBE8228"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.SI_36\(21),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37.Z_C3_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"96696996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.SI_36\(21),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.SI_152\(17));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_C3_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"DEED4884"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_515\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.SI_51\(6),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_C3_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"69969669"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_515\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.SI_51\(6),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.SI_167\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47.Z_C3_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"BE28"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_C1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_AXB1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47.Z_C3_LUT6_2_O5\: LUT3 
generic map(
  INIT => X"96"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.CIN\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_C1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46.Z_AXB1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47.Z_AXB2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_SN_M1_I_O2_LUT6_2_O6\: LUT2 
generic map(
  INIT => X"D"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_708\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_SN_M1_I_O2_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"000A000C"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.STKGEN_1_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"00002882"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7498_I\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SALSBS_1\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN12_GEN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN10_NOTPROP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.STKGEN_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.STKGEN_1_LUT6_2_O5\: LUT3 
generic map(
  INIT => X"9F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7498_I\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SALSBS_1\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN10_NOTPROP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.NOTPROP_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9.Z_C2_LUT6_2_O6\: LUT3 
generic map(
  INIT => X"E8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9.Z_C1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.SI_9\(48),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9.Z_C2_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"EDDE8448"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.CIN_1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.SI_9\(48),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10.Z_C2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33.Z_AXB2_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"6996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.SI_32\(25),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33.Z_AXB2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33.Z_AXB2_LUT6_2_O5\: LUT3 
generic map(
  INIT => X"E8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_C1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.SI_32\(25),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_AXB2_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"6996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.SI_28\(29),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_AXB2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29.Z_AXB2_LUT6_2_O5\: LUT3 
generic map(
  INIT => X"E8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28.Z_C1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.SI_28\(29),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28.Z_C2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_AC0_1_LUT6_2_O6\: LUT3 
generic map(
  INIT => X"48"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_C1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.SI_25\(32),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_AC0_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_AC0_1_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"6996"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.CIN_2\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.CIN\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_C1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.SI_25\(32),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26.Z_AXB2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN2_NOTDECODEDUNIMP_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"CFCFDFCF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(64),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(66),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(67),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.ENTRYPOINT\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN2_NOTDECODEDUNIMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN2_NOTDECODEDUNIMP_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"CFCFDFCF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(64),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(66),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(67),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.ENTRYPOINT\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN2_NOTDECODEDUNIMP_0_E\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_AC0_1_LUT6_2_O6\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_C1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_AXB1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_AC0_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_AC0_1_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"FEA8FAA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.CIN_1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_C1\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_AC0_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.SI_80\(33),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_AXB1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23.Z_C3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1_LUT6_2_O6[56]\: LUT4 
generic map(
  INIT => X"0028"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_M1_LUT6_2_O5[56]\: LUT5 
generic map(
  INIT => X"000C0CA0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(174),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7576_SN\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(57));
\GRLFPC20.COMB.UN1_R.I.EXC_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"0080"
)
port map (
  I0 => \GRLFPC20.R.I.EXC\(5),
  I1 => \GRLFPC20.R.I.V\,
  I2 => \GRLFPC20.COMB.V.I.EXEC_5\,
  I3 => \GRLFPC20.N_2000\,
  O => \GRLFPC20.N_2015\);
\GRLFPC20.COMB.UN1_R.I.EXC_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"55551555"
)
port map (
  I0 => \GRLFPC20.N_1295\,
  I1 => \GRLFPC20.R.I.EXC\(5),
  I2 => \GRLFPC20.R.I.V\,
  I3 => \GRLFPC20.COMB.V.I.EXEC_5\,
  I4 => \GRLFPC20.N_2000\,
  O => \GRLFPC20.N_1958\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_RNIRCGS3_O6\: LUT3 
generic map(
  INIT => X"80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO2_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_RNIRCGS3_O5\: LUT4 
generic map(
  INIT => X"8000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_3\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14.Z_AXBXC0_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"2DD2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(326),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(47),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.SI_15\(42));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14.Z_AXBXC0_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"D22D2DD2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(326),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(47),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.CIN_2\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15.Z_AXB1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41.Z_C1_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"F220"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(353),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(20),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.CIN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41.Z_C1_LUT6_2_O5\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(316),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_C1_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"F220"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(364),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(9),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_C1_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"2DD2D22D"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(364),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(9),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_499\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53.Z_AXB1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51.Z_C1_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"F220"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(363),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(10),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51.Z_C1_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"2DD2D22D"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(363),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(10),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_513\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52.Z_AXB1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37.Z_AXBXC0_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"2DD2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(349),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(24),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.SI_38\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37.Z_AXBXC0_LUT6_2_O5\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(360),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(13));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47.Z_AXBXC0_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"2DD2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(359),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(14),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.SI_48\(9));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47.Z_AXBXC0_LUT6_2_O5\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(352),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(21));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_AXB0_LUT6_2_O6\: LUT3 
generic map(
  INIT => X"D2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(342),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.CIN\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_AXB0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30.Z_AXB0_LUT6_2_O5\: LUT3 
generic map(
  INIT => X"D2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(337),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.CIN_3\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25.Z_AXB0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIL7DR_O6[314]\: LUT5 
generic map(
  INIT => X"F0660066"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(314),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(372),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(114),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN1_NOTPROP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIL7DR_O5[314]\: LUT5 
generic map(
  INIT => X"0F880088"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(314),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(372),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(114),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(8),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN3_GEN_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0_LUT6_2_O6[0]\: LUT4 
generic map(
  INIT => X"0F47"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(12),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0_LUT6_2_O5[0]\: LUT5 
generic map(
  INIT => X"3333505F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(12),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(56));
\GRLFPC20.FPI.OP2_LUT6_2_O6[32]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(0),
  I1 => rfo2_data2(0),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(32));
\GRLFPC20.FPI.OP2_LUT6_2_O5[32]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(1),
  I1 => rfo2_data2(1),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(33));
\GRLFPC20.FPI.OP2_LUT6_2_O6[35]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(3),
  I1 => rfo2_data2(3),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(35));
\GRLFPC20.FPI.OP2_LUT6_2_O5[35]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(4),
  I1 => rfo2_data2(4),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(36));
\GRLFPC20.FPI.OP2_LUT6_2_O6[37]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(5),
  I1 => rfo2_data2(5),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(37));
\GRLFPC20.FPI.OP2_LUT6_2_O5[37]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(6),
  I1 => rfo2_data2(6),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(38));
\GRLFPC20.FPI.OP2_LUT6_2_O6[39]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(7),
  I1 => rfo2_data2(7),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(39));
\GRLFPC20.FPI.OP2_LUT6_2_O5[39]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(12),
  I1 => rfo2_data2(12),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(44));
\GRLFPC20.FPI.OP2_LUT6_2_O6[40]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(8),
  I1 => rfo2_data2(8),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(40));
\GRLFPC20.FPI.OP2_LUT6_2_O5[40]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(9),
  I1 => rfo2_data2(9),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(41));
\GRLFPC20.FPI.OP2_LUT6_2_O6[42]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(10),
  I1 => rfo2_data2(10),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(42));
\GRLFPC20.FPI.OP2_LUT6_2_O5[42]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(11),
  I1 => rfo2_data2(11),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(43));
\GRLFPC20.FPI.OP2_LUT6_2_O6[45]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(13),
  I1 => rfo2_data2(13),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(45));
\GRLFPC20.FPI.OP2_LUT6_2_O5[45]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(14),
  I1 => rfo2_data2(14),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(46));
\GRLFPC20.FPI.OP2_LUT6_2_O6[47]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(15),
  I1 => rfo2_data2(15),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(47));
\GRLFPC20.FPI.OP2_LUT6_2_O5[47]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(16),
  I1 => rfo2_data2(16),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(48));
\GRLFPC20.FPI.OP2_LUT6_2_O6[49]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(17),
  I1 => rfo2_data2(17),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(49));
\GRLFPC20.FPI.OP2_LUT6_2_O5[49]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(18),
  I1 => rfo2_data2(18),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(50));
\GRLFPC20.FPI.OP2_LUT6_2_O6[51]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(19),
  I1 => rfo2_data2(19),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(51));
\GRLFPC20.FPI.OP2_LUT6_2_O5[51]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(22),
  I1 => rfo2_data2(22),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(54));
\GRLFPC20.FPI.OP2_LUT6_2_O6[52]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(20),
  I1 => rfo2_data2(20),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(52));
\GRLFPC20.FPI.OP2_LUT6_2_O5[52]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(21),
  I1 => rfo2_data2(21),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(53));
\GRLFPC20.FPI.OP2_LUT6_2_O6[55]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(23),
  I1 => rfo2_data2(23),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(55));
\GRLFPC20.FPI.OP2_LUT6_2_O5[55]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(24),
  I1 => rfo2_data2(24),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(56));
\GRLFPC20.FPI.OP2_LUT6_2_O6[57]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(25),
  I1 => rfo2_data2(25),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(57));
\GRLFPC20.FPI.OP2_LUT6_2_O5[57]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(26),
  I1 => rfo2_data2(26),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(58));
\GRLFPC20.FPI.OP2_LUT6_2_O6[59]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(27),
  I1 => rfo2_data2(27),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(59));
\GRLFPC20.FPI.OP2_LUT6_2_O5[59]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(28),
  I1 => rfo2_data2(28),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(60));
\GRLFPC20.FPI.OP2_LUT6_2_O6[61]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(29),
  I1 => rfo2_data2(29),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(61));
\GRLFPC20.FPI.OP2_LUT6_2_O5[61]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => rfo1_data2(30),
  I1 => rfo2_data2(30),
  I2 => \GRLFPC20.COMB.UN1_FPCI_4\,
  O => \GRLFPC20.FPI.OP2\(62));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0_LUT6_2_O6[9]\: LUT5 
generic map(
  INIT => X"3333550F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(243),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_95\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(48));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0_LUT6_2_O5[9]\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.LIB\(1));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_1_LUT6_2_O6[0]\: LUT4 
generic map(
  INIT => X"BF00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_29_REP1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8532\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_1_LUT6_2_O5[0]\: LUT4 
generic map(
  INIT => X"EC00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8533\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIPN2P1_1_O6[78]\: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_11378\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIPN2P1_1_O5[78]\: LUT4 
generic map(
  INIT => X"24A8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10016\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_18_LUT6_2_O6[29]\: LUT5 
generic map(
  INIT => X"00000008"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1283\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_18_LUT6_2_O5[29]\: LUT4 
generic map(
  INIT => X"A4E0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9596\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_9_1_LUT6_2_O6[57]\: LUT5 
generic map(
  INIT => X"00001300"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_9_1\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_9_1_LUT6_2_O5[57]\: LUT5 
generic map(
  INIT => X"14C000F0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9709\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1_0_LUT6_2_O6[4]\: LUT5 
generic map(
  INIT => X"00015555"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(246),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(248),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(249),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(247),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1_0\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1_0_LUT6_2_O5[4]\: LUT4 
generic map(
  INIT => X"007F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(248),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(249),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(247),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN4_NOTBINFNAN\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_1_LUT6_2_O6[3]\: LUT4 
generic map(
  INIT => X"CE00"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8535\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_1_LUT6_2_O5[3]\: LUT3 
generic map(
  INIT => X"E0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8534\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O2_LUT6_2_O6[32]\: LUT2 
generic map(
  INIT => X"9"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1561\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O2_LUT6_2_O5[32]\: LUT4 
generic map(
  INIT => X"4802"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10917\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_28_0_LUT6_2_O6[75]\: LUT5 
generic map(
  INIT => X"FFFFEEEF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(77),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(76),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(75),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14\(77),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_28_0\(75));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_28_0_LUT6_2_O5[75]\: LUT4 
generic map(
  INIT => X"1110"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(77),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(76),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(75),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CONDMUXMULXFF.UN5_NOTSQRTLFTCC\);
\GRLFPC20.UN1_FPOP7_0_O2_LUT6_2_O6\: LUT3 
generic map(
  INIT => X"62"
)
port map (
  I0 => cpi_d_inst(7),
  I1 => cpi_d_inst(9),
  I2 => cpi_d_inst(12),
  O => \GRLFPC20.N_3079\);
\GRLFPC20.UN1_FPOP7_0_O2_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"0C0E0000"
)
port map (
  I0 => cpi_d_inst(7),
  I1 => cpi_d_inst(9),
  I2 => cpi_d_inst(12),
  I3 => cpi_d_inst(8),
  I4 => cpi_d_inst(11),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_6_0_E\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_1_LUT6_2_O6[7]\: LUT4 
generic map(
  INIT => X"0800"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8539\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_1_LUT6_2_O5[7]\: LUT3 
generic map(
  INIT => X"08"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1137\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O2_1_LUT6_2_O6[0]\: LUT2 
generic map(
  INIT => X"9"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_759\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O2_1_LUT6_2_O5[0]\: LUT3 
generic map(
  INIT => X"81"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10724\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTAINFNAN_0_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"80000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(237),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(238),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(239),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(242),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(243),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTAINFNAN_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTAINFNAN_0_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"FFFE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(237),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(238),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(239),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(242),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_1_0\(5));
\GRLFPC20.COMB.V.A.LD_1_1_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"0B000000"
)
port map (
  I0 => cpi_d_inst(19),
  I1 => cpi_d_inst(20),
  I2 => cpi_d_inst(22),
  I3 => cpi_d_inst(30),
  I4 => cpi_d_inst(31),
  O => \GRLFPC20.COMB.V.A.LD_1_1\);
\GRLFPC20.COMB.V.A.LD_1_1_LUT6_2_O5\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => cpi_d_inst(30),
  I1 => cpi_d_inst(31),
  O => \GRLFPC20.N_878\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS_LUT6_2_O6[4]\: LUT4 
generic map(
  INIT => X"E020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(240),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS_LUT6_2_O5[4]\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1323\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIVNQN1_O6[107]\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_812_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIVNQN1_O5[107]\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_846_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.UN84_TEMP_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.UN84_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.UN84_TEMP_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.UN138_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.UN348_TEMP_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.UN348_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.UN348_TEMP_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.UN462_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_LUT6_2_O6[6]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_FAST\(10),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_LUT6_2_O5[6]\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.UN3_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_3_LUT6_2_O6[75]\: LUT3 
generic map(
  INIT => X"95"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(48),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(52),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8807\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_3_LUT6_2_O5[75]\: LUT4 
generic map(
  INIT => X"8000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(49),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(48),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(51),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(52),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_26_A0_1\(75));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI28FK1_O6[66]\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_811_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNI28FK1_O5[66]\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.UN195_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIO6162_O6[72]\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_803_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH_RNIO6162_O5[72]\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.UN213_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.UN18_TEMP_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.UN18_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.UN18_TEMP_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.UN111_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.UN36_TEMP_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.UN36_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.UN36_TEMP_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.UN66_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.UN180_TEMP_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.UN180_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.UN180_TEMP_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.UN255_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_I_M2_LUT6_2_O6[4]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_707\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_I_M2_LUT6_2_O5[4]\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.UN252_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O24_4_LUT6_2_O6[59]\: LUT2 
generic map(
  INIT => X"B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10734\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O24_4_LUT6_2_O5[59]\: LUT4 
generic map(
  INIT => X"04C4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_7_0\(48));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14_2_LUT6_2_O6[77]\: LUT3 
generic map(
  INIT => X"54"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(77),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(76),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(75),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14_2\(77));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_14_2_LUT6_2_O5[77]\: LUT4 
generic map(
  INIT => X"BBBF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(61),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(76),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(75),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.UN33_PCTRL_NEW_I_0\);
\GRLFPC20.COMB.FPDECODE.RDD5_0_A2_LUT6_2_O6\: LUT3 
generic map(
  INIT => X"01"
)
port map (
  I0 => cpi_d_inst(9),
  I1 => cpi_d_inst(12),
  I2 => cpi_d_inst(13),
  O => \GRLFPC20.N_3116\);
\GRLFPC20.COMB.FPDECODE.RDD5_0_A2_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"00000100"
)
port map (
  I0 => cpi_d_inst(9),
  I1 => cpi_d_inst(12),
  I2 => cpi_d_inst(13),
  I3 => cpi_d_inst(5),
  I4 => cpi_d_inst(6),
  O => \GRLFPC20.N_3127\);
\GRLFPC20.COMB.FPDECODE.FPOP2_0_A2_LUT6_2_O6\: LUT3 
generic map(
  INIT => X"20"
)
port map (
  I0 => cpi_d_inst(21),
  I1 => cpi_d_inst(22),
  I2 => cpi_d_inst(24),
  O => \GRLFPC20.N_3109\);
\GRLFPC20.COMB.FPDECODE.FPOP2_0_A2_LUT6_2_O5\: LUT3 
generic map(
  INIT => X"08"
)
port map (
  I0 => cpi_d_inst(24),
  I1 => cpi_d_inst(19),
  I2 => cpi_d_inst(20),
  O => \GRLFPC20.COMB.V.A.AFSR_1_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1_I_0_LUT6_2_O6[1]\: LUT3 
generic map(
  INIT => X"3B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(1),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_101\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1_I_0_LUT6_2_O5[1]\: LUT3 
generic map(
  INIT => X"3B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(2),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_99\);
\GRLFPC20.COMB.V.E.FPOP_1_LUT6_2_O6\: LUT3 
generic map(
  INIT => X"10"
)
port map (
  I0 => cpi_a_annul,
  I1 => cpi_a_trap,
  I2 => \GRLFPC20.R.A.FPOP\,
  O => \GRLFPC20.N_2931_1\);
\GRLFPC20.COMB.V.E.FPOP_1_LUT6_2_O5\: LUT3 
generic map(
  INIT => X"10"
)
port map (
  I0 => cpi_a_annul,
  I1 => cpi_a_trap,
  I2 => \GRLFPC20.R.A.AFSR\,
  O => \GRLFPC20.COMB.V.E.AFSR_1\);
\GRLFPC20.ANNULFPU_0_SQMUXA_LUT6_2_O6\: LUT3 
generic map(
  INIT => X"E0"
)
port map (
  I0 => cpi_m_annul,
  I1 => cpi_m_trap,
  I2 => \GRLFPC20.R.M.FPOP\,
  O => \GRLFPC20.N_1536\);
\GRLFPC20.ANNULFPU_0_SQMUXA_LUT6_2_O5\: LUT3 
generic map(
  INIT => X"10"
)
port map (
  I0 => cpi_m_annul,
  I1 => cpi_m_trap,
  I2 => \GRLFPC20.R.M.AFSR\,
  O => \GRLFPC20.COMB.V.X.AFSR_1\);
\GRLFPC20.ANNULFPU_0_SQMUXA_1_LUT6_2_O6\: LUT3 
generic map(
  INIT => X"E0"
)
port map (
  I0 => cpi_e_annul,
  I1 => cpi_e_trap,
  I2 => \GRLFPC20.R.E.FPOP\,
  O => \GRLFPC20.N_1537\);
\GRLFPC20.ANNULFPU_0_SQMUXA_1_LUT6_2_O5\: LUT3 
generic map(
  INIT => X"10"
)
port map (
  I0 => cpi_e_annul,
  I1 => cpi_e_trap,
  I2 => \GRLFPC20.R.E.AFSR\,
  O => \GRLFPC20.COMB.V.M.AFSR_1\);
\GRLFPC20.ANNULFPU_0_SQMUXA_2_LUT6_2_O6\: LUT3 
generic map(
  INIT => X"E0"
)
port map (
  I0 => cpi_a_annul,
  I1 => cpi_a_trap,
  I2 => \GRLFPC20.R.A.FPOP\,
  O => \GRLFPC20.N_1538\);
\GRLFPC20.ANNULFPU_0_SQMUXA_2_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"0000001F"
)
port map (
  I0 => cpi_a_annul,
  I1 => cpi_a_trap,
  I2 => \GRLFPC20.R.A.FPOP\,
  I3 => \GRLFPC20.N_1536\,
  I4 => \GRLFPC20.N_1537\,
  O => \GRLFPC20.N_1528\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_0_1_LUT6_2_O6[6]\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9861_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_0_1_LUT6_2_O5[6]\: LUT2 
generic map(
  INIT => X"9"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_722\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_4_1_0_A2_LUT6_2_O6[54]\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9797_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_4_1_0_A2_LUT6_2_O5[54]\: LUT3 
generic map(
  INIT => X"01"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2517_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN3_S_SQRT_1_LUT6_2_O6\: LUT3 
generic map(
  INIT => X"60"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9913_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN3_S_SQRT_1_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"40004080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A12_0_0\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_6_1_LUT6_2_O6[48]\: LUT3 
generic map(
  INIT => X"01"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10161_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_6_1_LUT6_2_O5[48]\: LUT3 
generic map(
  INIT => X"60"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2695\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNITR2P1_O6[79]\: LUT3 
generic map(
  INIT => X"02"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_7_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNITR2P1_O5[79]\: LUT3 
generic map(
  INIT => X"01"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A30_23_0\(58));
\GRLFPC20.R.I.EXC_RNIG21C4_O6[2]\: LUT5 
generic map(
  INIT => X"00007F00"
)
port map (
  I0 => cpi_dbg_enable,
  I1 => cpi_dbg_fsr,
  I2 => cpi_dbg_write,
  I3 => \GRLFPC20.R.I.EXC\(2),
  I4 => \GRLFPC20.COMB.V.FSR.AEXC_1_SN.N_7_MUX\,
  O => \GRLFPC20.R.I.EXC_M\(2));
\GRLFPC20.R.I.EXC_RNIG21C4_O5[2]\: LUT3 
generic map(
  INIT => X"80"
)
port map (
  I0 => cpi_dbg_enable,
  I1 => cpi_dbg_fsr,
  I2 => cpi_dbg_write,
  O => \GRLFPC20.N_1704\);
\GRLFPC20.COMB.UN1_R.I.V_LUT6_2_O6\: LUT3 
generic map(
  INIT => X"40"
)
port map (
  I0 => \GRLFPC20.R.I.EXEC\,
  I1 => \GRLFPC20.R.I.V\,
  I2 => \GRLFPC20.R.X.FPOP\,
  O => \GRLFPC20.COMB.UN1_R.I.V\);
\GRLFPC20.COMB.UN1_R.I.V_LUT6_2_O5\: LUT2 
generic map(
  INIT => X"1"
)
port map (
  I0 => \GRLFPC20.R.I.EXEC\,
  I1 => \GRLFPC20.R.X.FPOP\,
  O => \GRLFPC20.N_1502_1\);
\GRLFPC20.COMB.UN1_FPCI_0_LUT6_2_O6\: LUT3 
generic map(
  INIT => X"FE"
)
port map (
  I0 => cpi_flush,
  I1 => cpi_x_annul,
  I2 => cpi_x_trap,
  O => \GRLFPC20.N_1295\);
\GRLFPC20.COMB.UN1_FPCI_0_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"01000000"
)
port map (
  I0 => cpi_flush,
  I1 => cpi_x_annul,
  I2 => cpi_x_trap,
  I3 => holdn,
  I4 => \GRLFPC20.R.X.FPOP\,
  O => N_3710);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN3_NOTAZERODENORM_LUT6_2_O6\: LUT3 
generic map(
  INIT => X"FE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(235),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(234),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(236),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN3_NOTAZERODENORM\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN3_NOTAZERODENORM_LUT6_2_O5\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(235),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(236),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN8_NOTAINFNAN_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MAPMULXFF.UN4_UNIMPMAP_LUT6_2_O6\: LUT3 
generic map(
  INIT => X"F7"
)
port map (
  I0 => cpi_d_inst(9),
  I1 => cpi_d_inst(11),
  I2 => cpi_d_inst(12),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7596\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MAPMULXFF.UN4_UNIMPMAP_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"0800"
)
port map (
  I0 => cpi_d_inst(9),
  I1 => cpi_d_inst(11),
  I2 => cpi_d_inst(12),
  I3 => cpi_d_inst(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_5_0_E\(1));
\GRLFPC20.COMB.SEQERR.UN3_QNE_1_0_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"8000"
)
port map (
  I0 => cpi_d_inst(21),
  I1 => cpi_d_inst(24),
  I2 => cpi_d_inst(30),
  I3 => cpi_d_inst(31),
  O => \GRLFPC20.COMB.SEQERR.UN3_QNE_1_0\);
\GRLFPC20.COMB.SEQERR.UN3_QNE_1_0_LUT6_2_O5\: LUT3 
generic map(
  INIT => X"40"
)
port map (
  I0 => cpi_d_inst(30),
  I1 => cpi_d_inst(31),
  I2 => \GRLFPC20.N_940\,
  O => \GRLFPC20.N_925\);
\GRLFPC20.COMB.UN1_MEXC_1_0_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"135F"
)
port map (
  I0 => \GRLFPC20.R.I.EXC\(2),
  I1 => \GRLFPC20.R.I.EXC\(3),
  I2 => \GRLFPC20.R.FSR.TEM\(2),
  I3 => \GRLFPC20.R.FSR.TEM\(3),
  O => \GRLFPC20.COMB.UN1_MEXC_1_0\);
\GRLFPC20.COMB.UN1_MEXC_1_0_LUT6_2_O5\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.R.I.EXC\(3),
  I1 => \GRLFPC20.R.FSR.TEM\(3),
  O => \GRLFPC20.N_1309\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[60]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(53),
  I2 => N_3880,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9126\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[60]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(11),
  I2 => \GRLFPC20.FPO.FRAC\(13),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9084\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[92]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(21),
  I2 => \GRLFPC20.FPO.FRAC\(23),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9094\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[92]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(20),
  I2 => \GRLFPC20.FPO.FRAC\(22),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9093\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[70]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(43),
  I2 => \GRLFPC20.FPO.FRAC\(45),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9116\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[70]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(42),
  I2 => \GRLFPC20.FPO.FRAC\(44),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9115\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2_LUT6_2_O6[7]\: LUT3 
generic map(
  INIT => X"AC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(250),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(237),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8552\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2_LUT6_2_O5[7]\: LUT3 
generic map(
  INIT => X"AC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(251),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(238),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8551\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2_LUT6_2_O6[0]\: LUT3 
generic map(
  INIT => X"AC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(257),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8545\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2_LUT6_2_O5[0]\: LUT3 
generic map(
  INIT => X"AC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(252),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(239),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8550\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2_LUT6_2_O6[3]\: LUT3 
generic map(
  INIT => X"AC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(254),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(241),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8548\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2_LUT6_2_O5[3]\: LUT3 
generic map(
  INIT => X"AC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(253),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(240),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8549\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2_LUT6_2_O6[1]\: LUT3 
generic map(
  INIT => X"AC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(256),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(243),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8546\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2_LUT6_2_O5[1]\: LUT3 
generic map(
  INIT => X"AC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(255),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(242),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8547\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[77]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(36),
  I2 => \GRLFPC20.FPO.FRAC\(38),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9109\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[77]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(37),
  I2 => \GRLFPC20.FPO.FRAC\(39),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9110\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[107]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(6),
  I2 => \GRLFPC20.FPO.FRAC\(8),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9079\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[107]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(7),
  I2 => \GRLFPC20.FPO.FRAC\(9),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9080\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[87]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(26),
  I2 => \GRLFPC20.FPO.FRAC\(28),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9099\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[87]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(25),
  I2 => \GRLFPC20.FPO.FRAC\(27),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9098\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[83]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(30),
  I2 => \GRLFPC20.FPO.FRAC\(32),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9103\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[83]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(31),
  I2 => \GRLFPC20.FPO.FRAC\(33),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9104\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[79]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(34),
  I2 => \GRLFPC20.FPO.FRAC\(36),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9107\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[79]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(35),
  I2 => \GRLFPC20.FPO.FRAC\(37),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9108\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[81]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(32),
  I2 => \GRLFPC20.FPO.FRAC\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9105\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[81]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(33),
  I2 => \GRLFPC20.FPO.FRAC\(35),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9106\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[85]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(28),
  I2 => \GRLFPC20.FPO.FRAC\(30),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9101\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[85]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(29),
  I2 => \GRLFPC20.FPO.FRAC\(31),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9102\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[69]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(44),
  I2 => \GRLFPC20.FPO.FRAC\(46),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9117\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[69]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => N_3825,
  I2 => N_3827,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9073\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_LUT6_2_O6[2]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP1\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_LUT6_2_O5[2]\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.UN393_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[112]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => N_3826,
  I2 => \GRLFPC20.FPO.FRAC\(3),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9074\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[112]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => N_3827,
  I2 => \GRLFPC20.FPO.FRAC\(4),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9075\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[72]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(41),
  I2 => \GRLFPC20.FPO.FRAC\(43),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9114\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[72]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(3),
  I2 => \GRLFPC20.FPO.FRAC\(5),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9076\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[66]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(47),
  I2 => \GRLFPC20.FPO.FRAC\(49),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9120\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[66]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(8),
  I2 => \GRLFPC20.FPO.FRAC\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9081\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[104]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(9),
  I2 => \GRLFPC20.FPO.FRAC\(11),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9082\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[104]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(10),
  I2 => \GRLFPC20.FPO.FRAC\(12),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9083\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[101]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(12),
  I2 => \GRLFPC20.FPO.FRAC\(14),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9085\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[101]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(13),
  I2 => \GRLFPC20.FPO.FRAC\(15),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9086\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[97]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(16),
  I2 => \GRLFPC20.FPO.FRAC\(18),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9089\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[97]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(15),
  I2 => \GRLFPC20.FPO.FRAC\(17),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9088\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[62]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(51),
  I2 => \GRLFPC20.FPO.FRAC\(53),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9124\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[62]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(19),
  I2 => \GRLFPC20.FPO.FRAC\(21),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9092\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[91]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(22),
  I2 => \GRLFPC20.FPO.FRAC\(24),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9095\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[91]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(23),
  I2 => \GRLFPC20.FPO.FRAC\(25),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9096\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[89]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(24),
  I2 => \GRLFPC20.FPO.FRAC\(26),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9097\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[89]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(27),
  I2 => \GRLFPC20.FPO.FRAC\(29),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9100\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[74]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(39),
  I2 => \GRLFPC20.FPO.FRAC\(41),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9112\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[74]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(40),
  I2 => \GRLFPC20.FPO.FRAC\(42),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9113\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[67]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(46),
  I2 => \GRLFPC20.FPO.FRAC\(48),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9119\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[67]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(45),
  I2 => \GRLFPC20.FPO.FRAC\(47),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9118\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[65]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(48),
  I2 => \GRLFPC20.FPO.FRAC\(50),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9121\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[65]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(49),
  I2 => \GRLFPC20.FPO.FRAC\(51),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9122\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0_LUT6_2_O6[0]\: LUT3 
generic map(
  INIT => X"AC"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_10_REP2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0_LUT6_2_O5[0]\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.UN534_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2_LUT6_2_O6[8]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(236),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(249),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8553\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2_LUT6_2_O5[8]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(235),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(248),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8554\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[109]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(4),
  I2 => \GRLFPC20.FPO.FRAC\(6),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9077\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[109]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(5),
  I2 => \GRLFPC20.FPO.FRAC\(7),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9078\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[75]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(38),
  I2 => \GRLFPC20.FPO.FRAC\(40),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9111\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[75]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(14),
  I2 => \GRLFPC20.FPO.FRAC\(16),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9087\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O6[96]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(17),
  I2 => \GRLFPC20.FPO.FRAC\(19),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9090\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2_LUT6_2_O5[96]\: LUT3 
generic map(
  INIT => X"D8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
  I1 => \GRLFPC20.FPO.FRAC\(18),
  I2 => \GRLFPC20.FPO.FRAC\(20),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9091\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI4M721_1_O6[78]\: LUT2 
generic map(
  INIT => X"1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10948_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI4M721_1_O5[78]\: LUT2 
generic map(
  INIT => X"E"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_741\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_RNISJ7V2_O6[9]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1344\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_RNISJ7V2_O5[9]\: LUT4 
generic map(
  INIT => X"FF40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1006_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2502\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_FAST\(9));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A15_11_2_I_O2_LUT6_2_O6[18]\: LUT2 
generic map(
  INIT => X"B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_712\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A15_11_2_I_O2_LUT6_2_O5[18]\: LUT4 
generic map(
  INIT => X"FF40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1006_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2502\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(9));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.S_CMP_3_0_A2_I_O2_LUT6_2_O6\: LUT2 
generic map(
  INIT => X"E"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_717\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.S_CMP_3_0_A2_I_O2_LUT6_2_O5\: LUT2 
generic map(
  INIT => X"D"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_795\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_X2_LUT6_2_O6[60]\: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9296_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_X2_LUT6_2_O5[60]\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9670_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_6_2_LUT6_2_O6[25]\: LUT2 
generic map(
  INIT => X"1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9858_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_6_2_LUT6_2_O5[25]\: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_747_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_2_0_I_O2_LUT6_2_O6[57]\: LUT2 
generic map(
  INIT => X"B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10869\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_2_0_I_O2_LUT6_2_O5[57]\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9320_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_2_1_LUT6_2_O6[25]\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9973_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_2_1_LUT6_2_O5[25]\: LUT3 
generic map(
  INIT => X"10"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2724\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_17_1_LUT6_2_O6[32]\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1019_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_17_1_LUT6_2_O5[32]\: LUT2 
generic map(
  INIT => X"7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_52\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O26_5_I_A2_LUT6_2_O6[52]\: LUT2 
generic map(
  INIT => X"1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10207_I_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O26_5_I_A2_LUT6_2_O5[52]\: LUT4 
generic map(
  INIT => X"0020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9324_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_4_1_I_LUT6_2_O6[13]\: LUT2 
generic map(
  INIT => X"7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_125\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_4_1_I_LUT6_2_O5[13]\: LUT4 
generic map(
  INIT => X"0040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10891_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A12_8_1_LUT6_2_O6[0]\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9975_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A12_8_1_LUT6_2_O5[0]\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10824_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNITF821_O6[80]\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9389_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNITF821_O5[80]\: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12021_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI1V1P1_O6[78]\: LUT2 
generic map(
  INIT => X"7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_202\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI1V1P1_O5[78]\: LUT4 
generic map(
  INIT => X"4000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_8_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_X2_LUT6_2_O6[6]\: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9700_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_X2_LUT6_2_O5[6]\: LUT2 
generic map(
  INIT => X"7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_749\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_0_A2_I_O2_LUT6_2_O6[48]\: LUT2 
generic map(
  INIT => X"D"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_766\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_0_A2_I_O2_LUT6_2_O5[48]\: LUT5 
generic map(
  INIT => X"FFFF0040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_157_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_222\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1971\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1661\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI5N721_O6[79]\: LUT2 
generic map(
  INIT => X"7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_234\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI5N721_O5[79]\: LUT2 
generic map(
  INIT => X"7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_775\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_9_1_LUT6_2_O6[13]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9558_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_9_1_LUT6_2_O5[13]\: LUT2 
generic map(
  INIT => X"1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1048_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_14_1_LUT6_2_O6[6]\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9505_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_14_1_LUT6_2_O5[6]\: LUT2 
generic map(
  INIT => X"B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_16\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN6_S_11_2_0_A2_0_A2_0_A2_LUT6_2_O6\: LUT2 
generic map(
  INIT => X"1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9994_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN6_S_11_2_0_A2_0_A2_0_A2_LUT6_2_O5\: LUT2 
generic map(
  INIT => X"E"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_715\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_1_A2_RNI6K161_O6[37]\: LUT2 
generic map(
  INIT => X"7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_13\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_1_A2_RNI6K161_O5[37]\: LUT5 
generic map(
  INIT => X"FFFF0020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1580\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12131\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_969\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_1\(37));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI6O721_O6[79]\: LUT2 
generic map(
  INIT => X"7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9467\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI6O721_O5[79]\: LUT2 
generic map(
  INIT => X"7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_831\);
\GRLFPC20.COMB.RSDECODE.RS1V2_0_A2_0_LUT6_2_O6\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => cpi_d_inst(7),
  I1 => cpi_d_inst(8),
  O => \GRLFPC20.N_3123\);
\GRLFPC20.COMB.RSDECODE.RS1V2_0_A2_0_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"0040"
)
port map (
  I0 => cpi_d_inst(7),
  I1 => cpi_d_inst(9),
  I2 => cpi_d_inst(11),
  I3 => cpi_d_inst(12),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_4_0_E\(2));
\GRLFPC20.COMB.RDD_1.M4_E_I_A2_1_LUT6_2_O6\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => cpi_d_inst(5),
  I1 => cpi_d_inst(6),
  O => \GRLFPC20.N_3120\);
\GRLFPC20.COMB.RDD_1.M4_E_I_A2_1_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"FFFF44B0"
)
port map (
  I0 => cpi_d_inst(5),
  I1 => cpi_d_inst(6),
  I2 => \GRLFPC20.N_3082\,
  I3 => \GRLFPC20.N_3083_1\,
  I4 => \GRLFPC20.N_3084\,
  O => \GRLFPC20.N_3074\);
\GRLFPC20.COMB.RSDECODE.RS1V2_0_A2_LUT6_2_O6\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => cpi_d_inst(10),
  I1 => cpi_d_inst(11),
  O => \GRLFPC20.N_3117\);
\GRLFPC20.COMB.RSDECODE.RS1V2_0_A2_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"0400"
)
port map (
  I0 => cpi_d_inst(10),
  I1 => cpi_d_inst(11),
  I2 => cpi_d_inst(5),
  I3 => cpi_d_inst(6),
  O => \GRLFPC20.N_3128\);
\GRLFPC20.COMB.WRADDR_0_SQMUXA_LUT6_2_O6\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => \GRLFPC20.R.X.AFSR\,
  I1 => \GRLFPC20.R.X.LD\,
  O => \GRLFPC20.N_1475\);
\GRLFPC20.COMB.WRADDR_0_SQMUXA_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"E2F0F0F0"
)
port map (
  I0 => cpi_lddata(6),
  I1 => \GRLFPC20.N_1295\,
  I2 => \GRLFPC20.R.FSR.AEXC\(1),
  I3 => \GRLFPC20.R.X.AFSR\,
  I4 => \GRLFPC20.R.X.LD\,
  O => \GRLFPC20.COMB.V.FSR.AEXC_1_M0\(1));
\GRLFPC20.COMB.V.MK.BUSY_2_1_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"00080000"
)
port map (
  I0 => \GRLFPC20.R.MK.HOLDN2\,
  I1 => \GRLFPC20.R.MK.HOLDN1\,
  I2 => \GRLFPC20.R.MK.RST\,
  I3 => \GRLFPC20.R.MK.RST2\,
  I4 => \GRLFPC20.COMB.UN1_ANNULFPU\,
  O => \GRLFPC20.COMB.V.MK.BUSY_2_1\);
\GRLFPC20.COMB.V.MK.BUSY_2_1_LUT6_2_O5\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.R.MK.HOLDN2\,
  I1 => \GRLFPC20.R.MK.HOLDN1\,
  O => cpo_holdn);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16_LUT6_2_O6[45]\: LUT4 
generic map(
  INIT => X"04BF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(44),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(45),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(45));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16_LUT6_2_O5[45]\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(1),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1086\);
\GRLFPC20.COMB.V.E.STDATA2_LUT6_2_O6\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => cpi_a_cnt(0),
  I1 => cpi_a_cnt(1),
  O => \GRLFPC20.COMB.V.E.STDATA2\);
\GRLFPC20.COMB.V.E.STDATA2_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"F2D0"
)
port map (
  I0 => cpi_a_cnt(0),
  I1 => cpi_a_cnt(1),
  I2 => \GRLFPC20.R.I.INST\(6),
  I3 => \GRLFPC20.R.I.PC\(6),
  O => \GRLFPC20.N_2345\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A12_1_0_I_O2_LUT6_2_O6[0]\: LUT2 
generic map(
  INIT => X"7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_909\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A12_1_0_I_O2_LUT6_2_O5[0]\: LUT5 
generic map(
  INIT => X"44020000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9669_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9548\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_5_1_I_O2_LUT6_2_O6[32]\: LUT2 
generic map(
  INIT => X"7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_906\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_5_1_I_O2_LUT6_2_O5[32]\: LUT2 
generic map(
  INIT => X"7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12132\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_22_1_I_O2_LUT6_2_O6[19]\: LUT2 
generic map(
  INIT => X"7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_907\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_22_1_I_O2_LUT6_2_O5[19]\: LUT2 
generic map(
  INIT => X"1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9555_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIH9LD1_O6[78]\: LUT2 
generic map(
  INIT => X"7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_304\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIH9LD1_O5[78]\: LUT3 
generic map(
  INIT => X"80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9925_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIPN2P1_0_O6[78]\: LUT2 
generic map(
  INIT => X"B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_796\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIPN2P1_0_O5[78]\: LUT4 
generic map(
  INIT => X"0100"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_4_A2_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_9_LUT6_2_O6[35]\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9394_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_9_LUT6_2_O5[35]\: LUT2 
generic map(
  INIT => X"D"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_328\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_4_3_0_I_O2_LUT6_2_O6[25]\: LUT2 
generic map(
  INIT => X"D"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_783\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_4_3_0_I_O2_LUT6_2_O5[25]\: LUT2 
generic map(
  INIT => X"7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9666_1_I_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI4M721_0_O6[78]\: LUT2 
generic map(
  INIT => X"D"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_776\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI4M721_0_O5[78]\: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9887_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI4M721_O6[78]\: LUT2 
generic map(
  INIT => X"D"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_289\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI4M721_O5[78]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1229\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_X2_0_X2_LUT6_2_O6[19]\: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_768_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_X2_0_X2_LUT6_2_O5[19]\: LUT2 
generic map(
  INIT => X"E"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_205\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI1K821_O6[80]\: LUT2 
generic map(
  INIT => X"D"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_428\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI1K821_O5[80]\: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_767_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIMDKD1_O6[78]\: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_751_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIMDKD1_O5[78]\: LUT3 
generic map(
  INIT => X"40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9993\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_1_1_I_O2_LUT6_2_O6[25]\: LUT2 
generic map(
  INIT => X"7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9785_1_I_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_1_1_I_O2_LUT6_2_O5[25]\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9338_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIMK2P1_O6[78]\: LUT2 
generic map(
  INIT => X"E"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_732\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIMK2P1_O5[78]\: LUT4 
generic map(
  INIT => X"4000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A26_22_0\(60));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIPN2P1_O6[78]\: LUT2 
generic map(
  INIT => X"D"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_720\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIPN2P1_O5[78]\: LUT4 
generic map(
  INIT => X"00D0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A24_7_0\(59));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNID5LD1_O6[78]\: LUT2 
generic map(
  INIT => X"7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10410\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNID5LD1_O5[78]\: LUT3 
generic map(
  INIT => X"80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10441_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN3_S_SQRT_2_0_A2_0_A2_LUT6_2_O6\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9506_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN3_S_SQRT_2_0_A2_0_A2_LUT6_2_O5\: LUT2 
generic map(
  INIT => X"D"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_409\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O15_0_I_A2_I_LUT6_2_O6[18]\: LUT2 
generic map(
  INIT => X"E"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_406\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O15_0_I_A2_I_LUT6_2_O5[18]\: LUT5 
generic map(
  INIT => X"FFFFFF10"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2206\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2208\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19\(46));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_12_0_A2_I_LUT6_2_O6[62]\: LUT2 
generic map(
  INIT => X"B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_261\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_12_0_A2_I_LUT6_2_O5[62]\: LUT4 
generic map(
  INIT => X"0080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A30_4_1\(58));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_6_1_I_LUT6_2_O6[36]\: LUT2 
generic map(
  INIT => X"7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_76\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_6_1_I_LUT6_2_O5[36]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10025_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN7_S_14_2_I_LUT6_2_O6\: LUT2 
generic map(
  INIT => X"E"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_59\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN7_S_14_2_I_LUT6_2_O5\: LUT2 
generic map(
  INIT => X"1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9652_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O2_I_A2_I_LUT6_2_O6[47]\: LUT2 
generic map(
  INIT => X"E"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12195\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O2_I_A2_I_LUT6_2_O5[47]\: LUT3 
generic map(
  INIT => X"01"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9404_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_RNI1SP71_O6[28]\: LUT2 
generic map(
  INIT => X"1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9468_I_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_RNI1SP71_O5[28]\: LUT5 
generic map(
  INIT => X"FFFF2100"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2758\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2341\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_0\(28));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIQO2P1_O6[79]\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9508_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIQO2P1_O5[79]\: LUT4 
generic map(
  INIT => X"0800"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A30_14_0\(58));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_1_0_0_A2_LUT6_2_O6[32]\: LUT2 
generic map(
  INIT => X"1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9503_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_1_0_0_A2_LUT6_2_O5[32]\: LUT4 
generic map(
  INIT => X"0001"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_15_1\(36));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_2_2_LUT6_2_O6[48]\: LUT3 
generic map(
  INIT => X"20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10157_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_2_2_LUT6_2_O5[48]\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9563_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_1_1_0_A2_LUT6_2_O6[36]\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9738_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_1_1_0_A2_LUT6_2_O5[36]\: LUT2 
generic map(
  INIT => X"1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9850_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A15_2_2_0_A2_LUT6_2_O6[18]\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9601_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A15_2_2_0_A2_LUT6_2_O5[18]\: LUT2 
generic map(
  INIT => X"1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1149\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIF7LD1_O6[79]\: LUT2 
generic map(
  INIT => X"1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_291_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIF7LD1_O5[79]\: LUT3 
generic map(
  INIT => X"20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9666_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_5_1_0_A2_0_A2_LUT6_2_O6[13]\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9671_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_5_1_0_A2_0_A2_LUT6_2_O5[13]\: LUT2 
generic map(
  INIT => X"E"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_830\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6_LUT6_2_O6[41]\: LUT5 
generic map(
  INIT => X"003BC4FF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE\(1),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8214\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8216\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(41));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6_LUT6_2_O5[41]\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_187\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIH9LD1_0_O6[78]\: LUT2 
generic map(
  INIT => X"1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9972_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIH9LD1_0_O5[78]\: LUT3 
generic map(
  INIT => X"08"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10746_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI7O621_O6[78]\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9492_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI7O621_O5[78]\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9723_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI1J721_O6[78]\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_314_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI1J721_O5[78]\: LUT2 
generic map(
  INIT => X"1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9600_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_1_0_0_A2_LUT6_2_O6[61]\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10767_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_1_0_0_A2_LUT6_2_O5[61]\: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10592_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_5_2_0_A2_LUT6_2_O6[13]\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9790_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_5_2_0_A2_LUT6_2_O5[13]\: LUT4 
generic map(
  INIT => X"FF80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2707\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2336\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1654\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_0_2_0_A2_LUT6_2_O6[61]\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9969_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_0_2_0_A2_LUT6_2_O5[61]\: LUT2 
generic map(
  INIT => X"1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9576_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_O26_LUT6_2_O6[60]\: LUT2 
generic map(
  INIT => X"E"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10790\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_O26_LUT6_2_O5[60]\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9461_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_0_A2_0_A2_LUT6_2_O6[62]\: LUT3 
generic map(
  INIT => X"20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2583\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_0_A2_0_A2_LUT6_2_O5[62]\: LUT2 
generic map(
  INIT => X"B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9629\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O20_1_LUT6_2_O6[32]\: LUT2 
generic map(
  INIT => X"7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9828\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O20_1_LUT6_2_O5[32]\: LUT3 
generic map(
  INIT => X"32"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10236_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O2_LUT6_2_O6[36]\: LUT2 
generic map(
  INIT => X"B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10006\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O2_LUT6_2_O5[36]\: LUT3 
generic map(
  INIT => X"02"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2635\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O27_0_LUT6_2_O6[54]\: LUT2 
generic map(
  INIT => X"D"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10332\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O27_0_LUT6_2_O5[54]\: LUT4 
generic map(
  INIT => X"0040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1335\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_A2_12_LUT6_2_O6[31]\: LUT3 
generic map(
  INIT => X"20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9428\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_I_I_A2_12_LUT6_2_O5[31]\: LUT2 
generic map(
  INIT => X"B"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10576\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_4_1_LUT6_2_O6[61]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10888_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_4_1_LUT6_2_O5[61]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9610_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIF7LD1_O6[78]\: LUT3 
generic map(
  INIT => X"BF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_222\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIF7LD1_O5[78]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9968_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_4_2_LUT6_2_O6[32]\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9915_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_4_2_LUT6_2_O5[32]\: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10670_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_6_2_LUT6_2_O6[19]\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9657_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_6_2_LUT6_2_O5[19]\: LUT3 
generic map(
  INIT => X"09"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9390_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_2_1_LUT6_2_O6[13]\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9655_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_2_1_LUT6_2_O5[13]\: LUT3 
generic map(
  INIT => X"08"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2229_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_0_1_LUT6_2_O6[13]\: LUT2 
generic map(
  INIT => X"1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9549_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_0_1_LUT6_2_O5[13]\: LUT3 
generic map(
  INIT => X"04"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1272\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_5_1_LUT6_2_O6[6]\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1230\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_5_1_LUT6_2_O5[6]\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9969_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_9_1_LUT6_2_O6[6]\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9739_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_9_1_LUT6_2_O5[6]\: LUT4 
generic map(
  INIT => X"0200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_11_0\(19));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A12_7_1_LUT6_2_O6[0]\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9667_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A12_7_1_LUT6_2_O5[0]\: LUT5 
generic map(
  INIT => X"FFFFE000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9408_2\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2724\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9855\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_1_0\(7));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.S_CMP_2_LUT6_2_O6\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1132_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.S_CMP_2_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"0040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10694_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_X2_0_LUT6_2_O6[25]\: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9637_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_X2_0_LUT6_2_O5[25]\: LUT5 
generic map(
  INIT => X"FFFFFF40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_991_1\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3_0\(5),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_989\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_3\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_X2_LUT6_2_O6[52]\: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10584_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_X2_LUT6_2_O5[52]\: LUT5 
generic map(
  INIT => X"FFFF0070"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2635\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_742\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2230\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0\(15));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_X2_LUT6_2_O6[53]\: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9946_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_X2_LUT6_2_O5[53]\: LUT4 
generic map(
  INIT => X"40C0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_9_0\(55));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_X2_LUT6_2_O6[57]\: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10671_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_X2_LUT6_2_O5[57]\: LUT4 
generic map(
  INIT => X"0002"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2600\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O3_LUT6_2_O6[48]\: LUT2 
generic map(
  INIT => X"E"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10130\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O3_LUT6_2_O5[48]\: LUT4 
generic map(
  INIT => X"0008"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9857_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A15_5_1_LUT6_2_O6[18]\: LUT2 
generic map(
  INIT => X"8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9604_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A15_5_1_LUT6_2_O5[18]\: LUT4 
generic map(
  INIT => X"0010"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9669_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A15_6_1_LUT6_2_O6[18]\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9605_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A15_6_1_LUT6_2_O5[18]\: LUT4 
generic map(
  INIT => X"0020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10759_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_X2_LUT6_2_O6[25]\: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1536_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_X2_LUT6_2_O5[25]\: LUT3 
generic map(
  INIT => X"04"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2721\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_X2_LUT6_2_O6[34]\: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9366_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_X2_LUT6_2_O5[34]\: LUT4 
generic map(
  INIT => X"0080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2800\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_X2_1_LUT6_2_O6[52]\: LUT2 
generic map(
  INIT => X"6"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1553_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_X2_1_LUT6_2_O5[52]\: LUT3 
generic map(
  INIT => X"80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9916_1\);
\GRLFPC20.COMB.UN4_LOCK_RNISHUN_O6\: LUT2 
generic map(
  INIT => X"2"
)
port map (
  I0 => holdn,
  I1 => rst,
  O => N_3584);
\GRLFPC20.COMB.UN4_LOCK_RNISHUN_O5\: LUT3 
generic map(
  INIT => X"08"
)
port map (
  I0 => holdn,
  I1 => \GRLFPC20.N_1583\,
  I2 => \GRLFPC20.N_1317\,
  O => \GRLFPC20.RIN.MK.LDOP_0_E\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN10_S_MOV_0_LUT6_2_O6\: LUT2 
generic map(
  INIT => X"1"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9490_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN10_S_MOV_0_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"00000400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9328\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A26_16_0_LUT6_2_O6[60]\: LUT2 
generic map(
  INIT => X"4"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9911_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A26_16_0_LUT6_2_O5[60]\: LUT5 
generic map(
  INIT => X"C444C000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1011_1\,
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10891_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_5_0\(47));
\GRLFPC20.COMB.WREN1_11_IV_0_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"C4C0C4CC"
)
port map (
  I0 => cpi_x_inst(25),
  I1 => \GRLFPC20.N_2112\,
  I2 => \GRLFPC20.COMB.RDD_2\,
  I3 => \GRLFPC20.COMB.UN1_R.I.V\,
  I4 => \GRLFPC20.R.I.INST\(25),
  O => \GRLFPC20.COMB.WREN1_11_IV_0\);
\GRLFPC20.COMB.WREN1_11_IV_0_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"C8CCC8C0"
)
port map (
  I0 => cpi_x_inst(25),
  I1 => \GRLFPC20.N_2112\,
  I2 => \GRLFPC20.COMB.RDD_2\,
  I3 => \GRLFPC20.COMB.UN1_R.I.V\,
  I4 => \GRLFPC20.R.I.INST\(25),
  O => \GRLFPC20.COMB.WREN2_11_IV_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI0ICT1_O6[54]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(54),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_10\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI0ICT1_O5[54]\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(55),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_10\(5));
\GRLFPC20.FPI.START_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"00000008"
)
port map (
  I0 => holdn,
  I1 => \GRLFPC20.N_1583\,
  I2 => \GRLFPC20.R.MK.RST\,
  I3 => \GRLFPC20.R.MK.RST2\,
  I4 => \GRLFPC20.N_1317\,
  O => \GRLFPC20.FPI.START\);
\GRLFPC20.FPI.START_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"00000008"
)
port map (
  I0 => holdn,
  I1 => \GRLFPC20.N_1583\,
  I2 => \GRLFPC20.R.MK.RST\,
  I3 => \GRLFPC20.R.MK.RST2\,
  I4 => \GRLFPC20.N_1317\,
  O => \GRLFPC20.FPI.START_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_2_A2_1_A2_LUT6_2_O6[26]\: LUT4 
generic map(
  INIT => X"0800"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1192\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2380\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_2_A2_1_A2_LUT6_2_O5[26]\: LUT5 
generic map(
  INIT => X"80000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1192\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2214\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI0U1P1_O6[78]\: LUT4 
generic map(
  INIT => X"0004"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1192\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI0U1P1_O5[78]\: LUT4 
generic map(
  INIT => X"0100"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_2_0\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.UN537_TEMP_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.UN537_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.UN537_TEMP_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.UN543_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNID5LD1_0_O6[78]\: LUT3 
generic map(
  INIT => X"04"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1232\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNID5LD1_0_O5[78]\: LUT4 
generic map(
  INIT => X"0400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2608\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A24_18_1_LUT6_2_O6[59]\: LUT3 
generic map(
  INIT => X"20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10765_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A24_18_1_LUT6_2_O5[59]\: LUT4 
generic map(
  INIT => X"0200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1170\);
\GRLFPC20.V.FSR.NONSTD_0_SQMUXA_2_LUT6_2_O6\: LUT5 
generic map(
  INIT => X"01000000"
)
port map (
  I0 => cpi_flush,
  I1 => cpi_x_annul,
  I2 => cpi_x_trap,
  I3 => \GRLFPC20.R.X.AFSR\,
  I4 => \GRLFPC20.R.X.LD\,
  O => \GRLFPC20.N_1338\);
\GRLFPC20.V.FSR.NONSTD_0_SQMUXA_2_LUT6_2_O5\: LUT5 
generic map(
  INIT => X"00010000"
)
port map (
  I0 => cpi_flush,
  I1 => cpi_x_annul,
  I2 => cpi_x_trap,
  I3 => \GRLFPC20.R.X.AFSR\,
  I4 => \GRLFPC20.R.X.LD\,
  O => \GRLFPC20.N_1562\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_18_1_LUT6_2_O6[6]\: LUT3 
generic map(
  INIT => X"08"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9509_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_18_1_LUT6_2_O5[6]\: LUT3 
generic map(
  INIT => X"10"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A22_16_0\(53));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_17_2_LUT6_2_O6[55]\: LUT4 
generic map(
  INIT => X"0001"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10624_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_17_2_LUT6_2_O5[55]\: LUT4 
generic map(
  INIT => X"6401"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9957\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_5_A2_0_A2_I_LUT6_2_O6[51]\: LUT3 
generic map(
  INIT => X"F7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_398\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_5_A2_0_A2_I_LUT6_2_O5[51]\: LUT3 
generic map(
  INIT => X"20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_0\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.UN528_TEMP_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.UN528_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.UN528_TEMP_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.UN549_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_9_LUT6_2_O6[33]\: LUT3 
generic map(
  INIT => X"40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9941\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_9_LUT6_2_O5[33]\: LUT4 
generic map(
  INIT => X"0004"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9855_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_1_1_I_0_O2_LUT6_2_O6[48]\: LUT3 
generic map(
  INIT => X"7F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_135\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_1_1_I_0_O2_LUT6_2_O5[48]\: LUT3 
generic map(
  INIT => X"40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2590\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O27_5_LUT6_2_O6[33]\: LUT4 
generic map(
  INIT => X"F222"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9896\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O27_5_LUT6_2_O5[33]\: LUT4 
generic map(
  INIT => X"0080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9922_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_9_2_LUT6_2_O6[54]\: LUT4 
generic map(
  INIT => X"0020"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10383_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_9_2_LUT6_2_O5[54]\: LUT4 
generic map(
  INIT => X"0004"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_1_0\(36));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_15_2_LUT6_2_O6[32]\: LUT4 
generic map(
  INIT => X"2000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9863_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_15_2_LUT6_2_O5[32]\: LUT4 
generic map(
  INIT => X"BFFB"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_254\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_2_A2_0_A2_LUT6_2_O6[56]\: LUT4 
generic map(
  INIT => X"0100"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2594\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_2_A2_0_A2_LUT6_2_O5[56]\: LUT4 
generic map(
  INIT => X"2000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10246_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_6_1_LUT6_2_O6[32]\: LUT5 
generic map(
  INIT => X"000040C0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_6_1\(32));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_6_1_LUT6_2_O5[32]\: LUT5 
generic map(
  INIT => X"10504040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_6_0\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.UN639_TEMP_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.UN639_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.UN639_TEMP_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.UN546_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.UN555_TEMP_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.UN555_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.UN555_TEMP_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.UN633_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.UN531_TEMP_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.UN531_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.UN531_TEMP_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.UN552_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_16_LUT6_2_O6[29]\: LUT4 
generic map(
  INIT => X"0040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1169\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_16_LUT6_2_O5[29]\: LUT4 
generic map(
  INIT => X"0010"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10927_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.UN459_TEMP_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.UN459_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.UN459_TEMP_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"665A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.UN390_TEMP\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A30_4_0_LUT6_2_O6[58]\: LUT3 
generic map(
  INIT => X"45"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A30_4_0\(58));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A30_4_0_LUT6_2_O5[58]\: LUT3 
generic map(
  INIT => X"10"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9788_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_10_2_LUT6_2_O6[33]\: LUT3 
generic map(
  INIT => X"01"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9919_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_10_2_LUT6_2_O5[33]\: LUT4 
generic map(
  INIT => X"1000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_134_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_20_0_LUT6_2_O6[57]\: LUT4 
generic map(
  INIT => X"0001"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_20_0\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_20_0_LUT6_2_O5[57]\: LUT4 
generic map(
  INIT => X"0800"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1336\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_LUT6_2_O6[0]\: LUT3 
generic map(
  INIT => X"10"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2693\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_LUT6_2_O5[0]\: LUT3 
generic map(
  INIT => X"20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9408_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_14_1_LUT6_2_O6[27]\: LUT4 
generic map(
  INIT => X"0100"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9800_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_14_1_LUT6_2_O5[27]\: LUT4 
generic map(
  INIT => X"0001"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10626_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_1_I_0_O2_LUT6_2_O6[53]\: LUT3 
generic map(
  INIT => X"7F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12131\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_1_I_0_O2_LUT6_2_O5[53]\: LUT3 
generic map(
  INIT => X"10"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10752_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_3_2_LUT6_2_O6[49]\: LUT4 
generic map(
  INIT => X"0100"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2162_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_3_2_LUT6_2_O5[49]\: LUT4 
generic map(
  INIT => X"0400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10631_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O25_2_LUT6_2_O6[6]\: LUT3 
generic map(
  INIT => X"B8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9473\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O25_2_LUT6_2_O5[6]\: LUT5 
generic map(
  INIT => X"00000200"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2707\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_2_LUT6_2_O6[57]\: LUT3 
generic map(
  INIT => X"80"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10891_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_2_LUT6_2_O5[57]\: LUT5 
generic map(
  INIT => X"08000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2708\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_X2_LUT6_2_O6[54]\: LUT3 
generic map(
  INIT => X"95"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10343_I\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_X2_LUT6_2_O5[54]\: LUT3 
generic map(
  INIT => X"08"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9906_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A12_5_1_LUT6_2_O6[0]\: LUT3 
generic map(
  INIT => X"04"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1267\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A12_5_1_LUT6_2_O5[0]\: LUT3 
generic map(
  INIT => X"7F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_143\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNITT0D1_O6[5]\: LUT5 
generic map(
  INIT => X"00000020"
)
port map (
  I0 => rst,
  I1 => \GRLFPC20.R.MK.LDOP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(5),
  I3 => \GRLFPC20.R.MK.RST\,
  I4 => \GRLFPC20.R.MK.RST2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_N_6\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNITT0D1_O5[5]\: LUT3 
generic map(
  INIT => X"FD"
)
port map (
  I0 => rst,
  I1 => \GRLFPC20.R.MK.RST\,
  I2 => \GRLFPC20.R.MK.RST2\,
  O => \GRLFPC20.FPI.RST_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_14_4_LUT6_2_O6[32]\: LUT4 
generic map(
  INIT => X"0400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2701\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_14_4_LUT6_2_O5[32]\: LUT4 
generic map(
  INIT => X"0600"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_0_A2_0_A2_0\(51));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_3_0_LUT6_2_O6[55]\: LUT4 
generic map(
  INIT => X"0010"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10437_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_3_0_LUT6_2_O5[55]\: LUT5 
generic map(
  INIT => X"04000040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2505_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_24_2_LUT6_2_O6[57]\: LUT3 
generic map(
  INIT => X"08"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10629_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_24_2_LUT6_2_O5[57]\: LUT4 
generic map(
  INIT => X"0220"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_0\(15));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_5_LUT6_2_O6[57]\: LUT4 
generic map(
  INIT => X"0021"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10648\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_5_LUT6_2_O5[57]\: LUT4 
generic map(
  INIT => X"0004"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2697\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN1_ENTRYPOINT_0_LUT6_2_O6\: LUT3 
generic map(
  INIT => X"08"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_9_0\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN1_ENTRYPOINT_0_LUT6_2_O5\: LUT3 
generic map(
  INIT => X"08"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10696_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_5_4_LUT6_2_O6[61]\: LUT4 
generic map(
  INIT => X"0080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10693_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_5_4_LUT6_2_O5[61]\: LUT5 
generic map(
  INIT => X"00020000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A24_19_1\(59));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A2_5_LUT6_2_O6[60]\: LUT3 
generic map(
  INIT => X"20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10860\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A2_5_LUT6_2_O5[60]\: LUT3 
generic map(
  INIT => X"40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_7_0\(4));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_4_LUT6_2_O6[57]\: LUT4 
generic map(
  INIT => X"0C08"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10647\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_4_LUT6_2_O5[57]\: LUT4 
generic map(
  INIT => X"CC50"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10284\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_9_A2_0_A2_LUT6_2_O6[60]\: LUT3 
generic map(
  INIT => X"01"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2591\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_9_A2_0_A2_LUT6_2_O5[60]\: LUT3 
generic map(
  INIT => X"02"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10479\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_11_LUT6_2_O6[54]\: LUT3 
generic map(
  INIT => X"02"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10405\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_11_LUT6_2_O5[54]\: LUT4 
generic map(
  INIT => X"1000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1331\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_1_0_LUT6_2_O6[30]\: LUT4 
generic map(
  INIT => X"4000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2337_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_1_0_LUT6_2_O5[30]\: LUT3 
generic map(
  INIT => X"7F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9435\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_4_A2_0_A2_I_LUT6_2_O6[59]\: LUT3 
generic map(
  INIT => X"F7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_369\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_4_A2_0_A2_I_LUT6_2_O5[59]\: LUT3 
generic map(
  INIT => X"40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2797\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_13_LUT6_2_O6[24]\: LUT3 
generic map(
  INIT => X"08"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1175\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_13_LUT6_2_O5[24]\: LUT3 
generic map(
  INIT => X"F7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_411\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A30_12_LUT6_2_O6[58]\: LUT5 
generic map(
  INIT => X"00000100"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10690\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A30_12_LUT6_2_O5[58]\: LUT4 
generic map(
  INIT => X"0006"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1234\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_2_A2_0_A2_LUT6_2_O6[61]\: LUT3 
generic map(
  INIT => X"02"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_157_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_2_A2_0_A2_LUT6_2_O5[61]\: LUT3 
generic map(
  INIT => X"08"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A22_11_0\(53));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O2_3_A2_3_LUT6_2_O6[29]\: LUT4 
generic map(
  INIT => X"0001"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1333\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O2_3_A2_3_LUT6_2_O5[29]\: LUT5 
generic map(
  INIT => X"02000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10834\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O30_2_LUT6_2_O6[58]\: LUT3 
generic map(
  INIT => X"EF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10661\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O30_2_LUT6_2_O5[58]\: LUT5 
generic map(
  INIT => X"44000400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1562\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_1_I_LUT6_2_O6[47]\: LUT3 
generic map(
  INIT => X"7F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_595\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_1_I_LUT6_2_O5[47]\: LUT3 
generic map(
  INIT => X"01"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_0_0\(25));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_0_A2_0_A2_I_O2_LUT6_2_O6[61]\: LUT3 
generic map(
  INIT => X"F7"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_765\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_0_A2_0_A2_I_O2_LUT6_2_O5[61]\: LUT4 
generic map(
  INIT => X"0111"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_6081_A2_6_0\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_4_3_0_I_1_LUT6_2_O6[25]\: LUT3 
generic map(
  INIT => X"FD"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_12196_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_4_3_0_I_1_LUT6_2_O5[25]\: LUT3 
generic map(
  INIT => X"E0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9665_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI1V1P1_0_O6[78]\: LUT3 
generic map(
  INIT => X"10"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_999_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNI1V1P1_0_O5[78]\: LUT3 
generic map(
  INIT => X"01"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10943\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIUS2P1_O6[79]\: LUT3 
generic map(
  INIT => X"40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_990_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIUS2P1_O5[79]\: LUT3 
generic map(
  INIT => X"40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_0_0\(6));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_1_0_LUT6_2_O6[25]\: LUT4 
generic map(
  INIT => X"0080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_6095_A2_11_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_1_0_LUT6_2_O5[25]\: LUT5 
generic map(
  INIT => X"00004000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2758\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIML3P1_O6[80]\: LUT4 
generic map(
  INIT => X"0100"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_995_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_RNIML3P1_O5[80]\: LUT5 
generic map(
  INIT => X"08000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A24_10_1\(59));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15_0_A2_1_1_I_0_LUT6_2_O6[24]\: LUT3 
generic map(
  INIT => X"7F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_211\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_O15_0_A2_1_1_I_0_LUT6_2_O5[24]\: LUT3 
generic map(
  INIT => X"10"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2640\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O26_6_LUT6_2_O6[52]\: LUT3 
generic map(
  INIT => X"FE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10211\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O26_6_LUT6_2_O5[52]\: LUT3 
generic map(
  INIT => X"7F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_85\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A12_7_3_0_A2_0_A2_LUT6_2_O6[0]\: LUT3 
generic map(
  INIT => X"20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9453_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A12_7_3_0_A2_0_A2_LUT6_2_O5[0]\: LUT5 
generic map(
  INIT => X"00004000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2823\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_12_LUT6_2_O6[57]\: LUT3 
generic map(
  INIT => X"06"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10640\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_12_LUT6_2_O5[57]\: LUT3 
generic map(
  INIT => X"CE"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9642\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_11_LUT6_2_O6[57]\: LUT3 
generic map(
  INIT => X"D0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10654\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_11_LUT6_2_O5[57]\: LUT3 
generic map(
  INIT => X"21"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_0\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_2_A2_0_A2_LUT6_2_O6[59]\: LUT3 
generic map(
  INIT => X"10"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2584\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_2_A2_0_A2_LUT6_2_O5[59]\: LUT4 
generic map(
  INIT => X"00E0"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_6_0\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O20_3_LUT6_2_O6[32]\: LUT3 
generic map(
  INIT => X"F8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9840\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O20_3_LUT6_2_O5[32]\: LUT3 
generic map(
  INIT => X"B3"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10146\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_5_LUT6_2_O6[61]\: LUT3 
generic map(
  INIT => X"20"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2645\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_5_LUT6_2_O5[61]\: LUT3 
generic map(
  INIT => X"10"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_2_0\(5));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_6_1_LUT6_2_O6[11]\: LUT3 
generic map(
  INIT => X"C8"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9321_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_6_1_LUT6_2_O5[11]\: LUT5 
generic map(
  INIT => X"80000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1347\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_6_0_A2_I_O2_LUT6_2_O6[58]\: LUT3 
generic map(
  INIT => X"FB"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_921\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_6_0_A2_I_O2_LUT6_2_O5[58]\: LUT3 
generic map(
  INIT => X"42"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1580\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_7_LUT6_2_O6[61]\: LUT3 
generic map(
  INIT => X"04"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2669\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_7_LUT6_2_O5[61]\: LUT4 
generic map(
  INIT => X"0201"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_2_A2_0_A2_0\(51));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_0_LUT6_2_O6[61]\: LUT3 
generic map(
  INIT => X"02"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10895\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_0_LUT6_2_O5[61]\: LUT5 
generic map(
  INIT => X"00000080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1282\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A26_14_2_LUT6_2_O6[60]\: LUT3 
generic map(
  INIT => X"40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10087_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A26_14_2_LUT6_2_O5[60]\: LUT3 
generic map(
  INIT => X"40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_8_0\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_2_A2_1_A2_0_LUT6_2_O6[26]\: LUT5 
generic map(
  INIT => X"00000040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1342\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_2_A2_1_A2_0_LUT6_2_O5[26]\: LUT3 
generic map(
  INIT => X"08"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A12_0\(0));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_1_A2_0_A2_LUT6_2_O6[56]\: LUT4 
generic map(
  INIT => X"0002"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2606\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_1_A2_0_A2_LUT6_2_O5[56]\: LUT4 
generic map(
  INIT => X"4000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1011_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_1_1_LUT6_2_O6[36]\: LUT5 
generic map(
  INIT => X"00080000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_1_1\(36));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A15_1_1_LUT6_2_O5[36]\: LUT5 
generic map(
  INIT => X"00000450"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10948\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_7_1_LUT6_2_O6[25]\: LUT4 
generic map(
  INIT => X"2000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_7_1\(25));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_7_1_LUT6_2_O5[25]\: LUT4 
generic map(
  INIT => X"0504"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2454_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_6_0_LUT6_2_O6[57]\: LUT4 
generic map(
  INIT => X"1040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_6_0\(57));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A29_6_0_LUT6_2_O5[57]\: LUT4 
generic map(
  INIT => X"4000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_9_0\(25));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_6_I_O2_LUT6_2_O6[29]\: LUT3 
generic map(
  INIT => X"FD"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_742\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_6_I_O2_LUT6_2_O5[29]\: LUT4 
generic map(
  INIT => X"0010"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2605\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_11_1_LUT6_2_O6[13]\: LUT3 
generic map(
  INIT => X"10"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9560_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A19_11_1_LUT6_2_O5[13]\: LUT3 
generic map(
  INIT => X"10"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_23_0\(47));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_7_2_LUT6_2_O6[6]\: LUT4 
generic map(
  INIT => X"0800"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9664_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_7_2_LUT6_2_O5[6]\: LUT5 
generic map(
  INIT => X"00000080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_22_0\(54));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_11_0_LUT6_2_O6[52]\: LUT3 
generic map(
  INIT => X"8A"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_11_0\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_11_0_LUT6_2_O5[52]\: LUT5 
generic map(
  INIT => X"00304400"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => N_3154_TZ);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_10_1_LUT6_2_O6[61]\: LUT4 
generic map(
  INIT => X"0800"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_10_1\(61));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A13_10_1_LUT6_2_O5[61]\: LUT5 
generic map(
  INIT => X"00008000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_742\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1047\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_7_0_LUT6_2_O6[52]\: LUT4 
generic map(
  INIT => X"0060"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_7_0\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_7_0_LUT6_2_O5[52]\: LUT4 
generic map(
  INIT => X"0015"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_0_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A24_14_0_LUT6_2_O6[59]\: LUT4 
generic map(
  INIT => X"0080"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A26_16_0\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A24_14_0_LUT6_2_O5[59]\: LUT4 
generic map(
  INIT => X"0102"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A20_5_0\(48));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_17_0_LUT6_2_O6[33]\: LUT4 
generic map(
  INIT => X"4000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_17_0\(11));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A27_17_0_LUT6_2_O5[33]\: LUT5 
generic map(
  INIT => X"00004000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2706\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_10_0_LUT6_2_O6[6]\: LUT4 
generic map(
  INIT => X"0800"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9748\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A25_10_0_LUT6_2_O5[6]\: LUT5 
generic map(
  INIT => X"00080000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1002_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_5_0_LUT6_2_O6[35]\: LUT3 
generic map(
  INIT => X"10"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10223_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_A2_5_0_LUT6_2_O5[35]\: LUT5 
generic map(
  INIT => X"02000000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  I4 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2724\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_981\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_4_LUT6_2_O6[61]\: LUT4 
generic map(
  INIT => X"4000"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_2630\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_A2_4_LUT6_2_O5[61]\: LUT3 
generic map(
  INIT => X"40"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9577\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O2_4_LUT6_2_O6[29]\: LUT4 
generic map(
  INIT => X"0016"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_777\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_O2_4_LUT6_2_O5[29]\: LUT3 
generic map(
  INIT => X"08"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_10293_1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_1_1_LUT6_2_O6[11]\: LUT3 
generic map(
  INIT => X"01"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_9330_2\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_I_A27_1_1_LUT6_2_O5[11]\: LUT4 
generic map(
  INIT => X"0040"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1171\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4.Z_C1_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"F220"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(316),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4.Z_C1_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"2DD2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(316),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_5\(52));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54.Z_AXBXC0_LUT6_2_O6\: LUT4 
generic map(
  INIT => X"2DD2"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(366),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.SI_55\(2));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54.Z_AXBXC0_LUT6_2_O5\: LUT4 
generic map(
  INIT => X"F220"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(366),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(7),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.CIN_2\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54.Z_C1\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16_LUT6_2_O6[24]\: LUT4 
generic map(
  INIT => X"0B4F"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(24),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(23),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(24));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16_LUT6_2_O5[24]\: LUT4 
generic map(
  INIT => X"04BF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(24),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(25),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(25));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16_LUT6_2_O6[20]\: LUT4 
generic map(
  INIT => X"40FB"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(18),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(20),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(20));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16_LUT6_2_O5[20]\: LUT4 
generic map(
  INIT => X"04BF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(20),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(21),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(21));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16_LUT6_2_O6[23]\: LUT4 
generic map(
  INIT => X"04BF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(22),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(23),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(23));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16_LUT6_2_O5[23]\: LUT4 
generic map(
  INIT => X"04BF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(21),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(22),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(22));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16_LUT6_2_O6[44]\: LUT4 
generic map(
  INIT => X"04BF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(43),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(44),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(44));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16_LUT6_2_O5[44]\: LUT4 
generic map(
  INIT => X"04BF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8216\,
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(43),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(43));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16_LUT6_2_O6[12]\: LUT4 
generic map(
  INIT => X"40FB"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(10),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(12),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(12));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16_LUT6_2_O5[12]\: LUT4 
generic map(
  INIT => X"04BF"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(12),
  I3 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(13),
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(13));
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_39_U_N_3L3_LUT6_2_O6\: LUT3 
generic map(
  INIT => X"31"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(22),
  I1 => \GRLFPC20.FPI.LDOP\,
  I2 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.NOTABORTWB\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_39_U_N_3_3\);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_39_U_N_3L3_LUT6_2_O5\: LUT3 
generic map(
  INIT => X"CA"
)
port map (
  I0 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_8782\,
  I1 => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41\(253),
  I2 => \GRLFPC20.FPI.LDOP\,
  O => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(253));
cpo_exc <= CPO_EXC_1;
cpo_cc(0) <= NN_1;
cpo_cc(1) <= CPO_CC_3;
rfi1_rd1addr(0) <= RFI2_RD1ADDR_16;
rfi1_rd1addr(1) <= RFI2_RD1ADDR_17;
rfi1_rd1addr(2) <= RFI2_RD1ADDR_18;
rfi1_rd1addr(3) <= RFI2_RD1ADDR_19;
rfi1_rd2addr(0) <= RFI2_RD2ADDR_20;
rfi1_rd2addr(1) <= RFI2_RD2ADDR_21;
rfi1_rd2addr(2) <= RFI2_RD2ADDR_22;
rfi1_rd2addr(3) <= RFI2_RD2ADDR_23;
rfi1_wraddr(0) <= RFI2_WRADDR_24;
rfi1_wraddr(1) <= RFI2_WRADDR_25;
rfi1_wraddr(2) <= RFI2_WRADDR_26;
rfi1_wraddr(3) <= RFI2_WRADDR_27;
rfi2_rd1addr(0) <= RFI2_RD1ADDR_16;
rfi2_rd1addr(1) <= RFI2_RD1ADDR_17;
rfi2_rd1addr(2) <= RFI2_RD1ADDR_18;
rfi2_rd1addr(3) <= RFI2_RD1ADDR_19;
rfi2_rd2addr(0) <= RFI2_RD2ADDR_20;
rfi2_rd2addr(1) <= RFI2_RD2ADDR_21;
rfi2_rd2addr(2) <= RFI2_RD2ADDR_22;
rfi2_rd2addr(3) <= RFI2_RD2ADDR_23;
rfi2_wraddr(0) <= RFI2_WRADDR_24;
rfi2_wraddr(1) <= RFI2_WRADDR_25;
rfi2_wraddr(2) <= RFI2_WRADDR_26;
rfi2_wraddr(3) <= RFI2_WRADDR_27;
end beh;

