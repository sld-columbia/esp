../ariane/riscv_plic_wrap.sv