-- GRCAN 2.0 interface
  constant CFG_GRCAN       : integer := CONFIG_GRCAN_ENABLE;
  constant CFG_GRCANIRQ    : integer := CONFIG_GRCANIRQ;
  constant CFG_GRCANSINGLE : integer := CONFIG_GRCANSINGLE;

