../vortex/hw/rtl/tex_unit/VX_tex_define.vh