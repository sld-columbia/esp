
package version is
  constant grlib_version : integer := 1500;
  constant grlib_build : integer := 4164;
end;
