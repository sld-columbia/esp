../vortex/hw/rtl/VX_gpu_types.vh