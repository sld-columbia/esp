// ${ARIANE}/include/ariane_axi_pkg.sv requires these params defined here

package ariane_soc;

    localparam IdWidth = 4;
    localparam IdWidthSlave = IdWidth;

endpackage
