../vortex/hw/dpi/float_dpi.vh