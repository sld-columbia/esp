-- UART 1
  constant CFG_UART1_ENABLE : integer := CONFIG_UART1_ENABLE;
  constant CFG_UART1_FIFO   : integer := CFG_UA1_FIFO;
  constant CFG_UART1_IRQ : integer := CONFIG_UA1_IRQ;

